module os_64bit ( z0, z1, z2, y );
input [62:0] z0;
input [62:0] z1;
input [62:0] z2;
output [62:0] y;
wire [62:0] _y;
wire [62:0] _z0;
wire [62:0] _z1;
wire [62:0] _z2;
wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;
assign _z0 = z0;
assign _z1 = z1;
assign _z2 = z2;
assign y = _y;
XOR2UD1BWP30P140 U0 ( .A1( _z2[0] ), .A2( _z0[32] ), .Z( n0 ) );
XOR2UD1BWP30P140 U1 ( .A1( _z2[1] ), .A2( _z0[33] ), .Z( n1 ) );
XOR2UD1BWP30P140 U2 ( .A1( _z2[2] ), .A2( _z0[34] ), .Z( n2 ) );
XOR2UD1BWP30P140 U3 ( .A1( _z2[3] ), .A2( _z0[35] ), .Z( n3 ) );
XOR2UD1BWP30P140 U4 ( .A1( _z2[4] ), .A2( _z0[36] ), .Z( n4 ) );
XOR2UD1BWP30P140 U5 ( .A1( _z2[5] ), .A2( _z0[37] ), .Z( n5 ) );
XOR2UD1BWP30P140 U6 ( .A1( _z2[6] ), .A2( _z0[38] ), .Z( n6 ) );
XOR2UD1BWP30P140 U7 ( .A1( _z2[7] ), .A2( _z0[39] ), .Z( n7 ) );
XOR2UD1BWP30P140 U8 ( .A1( _z2[8] ), .A2( _z0[40] ), .Z( n8 ) );
XOR2UD1BWP30P140 U9 ( .A1( _z2[9] ), .A2( _z0[41] ), .Z( n9 ) );
XOR2UD1BWP30P140 U10 ( .A1( _z2[10] ), .A2( _z0[42] ), .Z( n10 ) );
XOR2UD1BWP30P140 U11 ( .A1( _z2[11] ), .A2( _z0[43] ), .Z( n11 ) );
XOR2UD1BWP30P140 U12 ( .A1( _z2[12] ), .A2( _z0[44] ), .Z( n12 ) );
XOR2UD1BWP30P140 U13 ( .A1( _z2[13] ), .A2( _z0[45] ), .Z( n13 ) );
XOR2UD1BWP30P140 U14 ( .A1( _z2[14] ), .A2( _z0[46] ), .Z( n14 ) );
XOR2UD1BWP30P140 U15 ( .A1( _z2[15] ), .A2( _z0[47] ), .Z( n15 ) );
XOR2UD1BWP30P140 U16 ( .A1( _z2[16] ), .A2( _z0[48] ), .Z( n16 ) );
XOR2UD1BWP30P140 U17 ( .A1( _z2[17] ), .A2( _z0[49] ), .Z( n17 ) );
XOR2UD1BWP30P140 U18 ( .A1( _z2[18] ), .A2( _z0[50] ), .Z( n18 ) );
XOR2UD1BWP30P140 U19 ( .A1( _z2[19] ), .A2( _z0[51] ), .Z( n19 ) );
XOR2UD1BWP30P140 U20 ( .A1( _z2[20] ), .A2( _z0[52] ), .Z( n20 ) );
XOR2UD1BWP30P140 U21 ( .A1( _z2[21] ), .A2( _z0[53] ), .Z( n21 ) );
XOR2UD1BWP30P140 U22 ( .A1( _z2[22] ), .A2( _z0[54] ), .Z( n22 ) );
XOR2UD1BWP30P140 U23 ( .A1( _z2[23] ), .A2( _z0[55] ), .Z( n23 ) );
XOR2UD1BWP30P140 U24 ( .A1( _z2[24] ), .A2( _z0[56] ), .Z( n24 ) );
XOR2UD1BWP30P140 U25 ( .A1( _z2[25] ), .A2( _z0[57] ), .Z( n25 ) );
XOR2UD1BWP30P140 U26 ( .A1( _z2[26] ), .A2( _z0[58] ), .Z( n26 ) );
XOR2UD1BWP30P140 U27 ( .A1( _z2[27] ), .A2( _z0[59] ), .Z( n27 ) );
XOR2UD1BWP30P140 U28 ( .A1( _z2[28] ), .A2( _z0[60] ), .Z( n28 ) );
XOR2UD1BWP30P140 U29 ( .A1( _z2[29] ), .A2( _z0[61] ), .Z( n29 ) );
XOR2UD1BWP30P140 U30 ( .A1( _z2[30] ), .A2( _z0[62] ), .Z( n30 ) );
XOR3UD1BWP30P140 U31 ( .A1( _z1[0] ), .A2( _z0[0] ), .A3( n0 ), .Z( _y[0] ) );
XOR3UD1BWP30P140 U32 ( .A1( _z1[1] ), .A2( _z0[1] ), .A3( n1 ), .Z( _y[1] ) );
XOR3UD1BWP30P140 U33 ( .A1( _z1[2] ), .A2( _z0[2] ), .A3( n2 ), .Z( _y[2] ) );
XOR3UD1BWP30P140 U34 ( .A1( _z1[3] ), .A2( _z0[3] ), .A3( n3 ), .Z( _y[3] ) );
XOR3UD1BWP30P140 U35 ( .A1( _z1[4] ), .A2( _z0[4] ), .A3( n4 ), .Z( _y[4] ) );
XOR3UD1BWP30P140 U36 ( .A1( _z1[5] ), .A2( _z0[5] ), .A3( n5 ), .Z( _y[5] ) );
XOR3UD1BWP30P140 U37 ( .A1( _z1[6] ), .A2( _z0[6] ), .A3( n6 ), .Z( _y[6] ) );
XOR3UD1BWP30P140 U38 ( .A1( _z1[7] ), .A2( _z0[7] ), .A3( n7 ), .Z( _y[7] ) );
XOR3UD1BWP30P140 U39 ( .A1( _z1[8] ), .A2( _z0[8] ), .A3( n8 ), .Z( _y[8] ) );
XOR3UD1BWP30P140 U40 ( .A1( _z1[9] ), .A2( _z0[9] ), .A3( n9 ), .Z( _y[9] ) );
XOR3UD1BWP30P140 U41 ( .A1( _z1[10] ), .A2( _z0[10] ), .A3( n10 ), .Z( _y[10] ) );
XOR3UD1BWP30P140 U42 ( .A1( _z1[11] ), .A2( _z0[11] ), .A3( n11 ), .Z( _y[11] ) );
XOR3UD1BWP30P140 U43 ( .A1( _z1[12] ), .A2( _z0[12] ), .A3( n12 ), .Z( _y[12] ) );
XOR3UD1BWP30P140 U44 ( .A1( _z1[13] ), .A2( _z0[13] ), .A3( n13 ), .Z( _y[13] ) );
XOR3UD1BWP30P140 U45 ( .A1( _z1[14] ), .A2( _z0[14] ), .A3( n14 ), .Z( _y[14] ) );
XOR3UD1BWP30P140 U46 ( .A1( _z1[15] ), .A2( _z0[15] ), .A3( n15 ), .Z( _y[15] ) );
XOR3UD1BWP30P140 U47 ( .A1( _z1[16] ), .A2( _z0[16] ), .A3( n16 ), .Z( _y[16] ) );
XOR3UD1BWP30P140 U48 ( .A1( _z1[17] ), .A2( _z0[17] ), .A3( n17 ), .Z( _y[17] ) );
XOR3UD1BWP30P140 U49 ( .A1( _z1[18] ), .A2( _z0[18] ), .A3( n18 ), .Z( _y[18] ) );
XOR3UD1BWP30P140 U50 ( .A1( _z1[19] ), .A2( _z0[19] ), .A3( n19 ), .Z( _y[19] ) );
XOR3UD1BWP30P140 U51 ( .A1( _z1[20] ), .A2( _z0[20] ), .A3( n20 ), .Z( _y[20] ) );
XOR3UD1BWP30P140 U52 ( .A1( _z1[21] ), .A2( _z0[21] ), .A3( n21 ), .Z( _y[21] ) );
XOR3UD1BWP30P140 U53 ( .A1( _z1[22] ), .A2( _z0[22] ), .A3( n22 ), .Z( _y[22] ) );
XOR3UD1BWP30P140 U54 ( .A1( _z1[23] ), .A2( _z0[23] ), .A3( n23 ), .Z( _y[23] ) );
XOR3UD1BWP30P140 U55 ( .A1( _z1[24] ), .A2( _z0[24] ), .A3( n24 ), .Z( _y[24] ) );
XOR3UD1BWP30P140 U56 ( .A1( _z1[25] ), .A2( _z0[25] ), .A3( n25 ), .Z( _y[25] ) );
XOR3UD1BWP30P140 U57 ( .A1( _z1[26] ), .A2( _z0[26] ), .A3( n26 ), .Z( _y[26] ) );
XOR3UD1BWP30P140 U58 ( .A1( _z1[27] ), .A2( _z0[27] ), .A3( n27 ), .Z( _y[27] ) );
XOR3UD1BWP30P140 U59 ( .A1( _z1[28] ), .A2( _z0[28] ), .A3( n28 ), .Z( _y[28] ) );
XOR3UD1BWP30P140 U60 ( .A1( _z1[29] ), .A2( _z0[29] ), .A3( n29 ), .Z( _y[29] ) );
XOR3UD1BWP30P140 U61 ( .A1( _z1[30] ), .A2( _z0[30] ), .A3( n30 ), .Z( _y[30] ) );
XOR3UD1BWP30P140 U62 ( .A1( _z2[31] ), .A2( _z1[31] ), .A3( _z0[31] ), .Z( _y[31] ) );
XOR3UD1BWP30P140 U63 ( .A1( _z1[32] ), .A2( _z2[32] ), .A3( n0 ), .Z( _y[32] ) );
XOR3UD1BWP30P140 U64 ( .A1( _z1[33] ), .A2( _z2[33] ), .A3( n1 ), .Z( _y[33] ) );
XOR3UD1BWP30P140 U65 ( .A1( _z1[34] ), .A2( _z2[34] ), .A3( n2 ), .Z( _y[34] ) );
XOR3UD1BWP30P140 U66 ( .A1( _z1[35] ), .A2( _z2[35] ), .A3( n3 ), .Z( _y[35] ) );
XOR3UD1BWP30P140 U67 ( .A1( _z1[36] ), .A2( _z2[36] ), .A3( n4 ), .Z( _y[36] ) );
XOR3UD1BWP30P140 U68 ( .A1( _z1[37] ), .A2( _z2[37] ), .A3( n5 ), .Z( _y[37] ) );
XOR3UD1BWP30P140 U69 ( .A1( _z1[38] ), .A2( _z2[38] ), .A3( n6 ), .Z( _y[38] ) );
XOR3UD1BWP30P140 U70 ( .A1( _z1[39] ), .A2( _z2[39] ), .A3( n7 ), .Z( _y[39] ) );
XOR3UD1BWP30P140 U71 ( .A1( _z1[40] ), .A2( _z2[40] ), .A3( n8 ), .Z( _y[40] ) );
XOR3UD1BWP30P140 U72 ( .A1( _z1[41] ), .A2( _z2[41] ), .A3( n9 ), .Z( _y[41] ) );
XOR3UD1BWP30P140 U73 ( .A1( _z1[42] ), .A2( _z2[42] ), .A3( n10 ), .Z( _y[42] ) );
XOR3UD1BWP30P140 U74 ( .A1( _z1[43] ), .A2( _z2[43] ), .A3( n11 ), .Z( _y[43] ) );
XOR3UD1BWP30P140 U75 ( .A1( _z1[44] ), .A2( _z2[44] ), .A3( n12 ), .Z( _y[44] ) );
XOR3UD1BWP30P140 U76 ( .A1( _z1[45] ), .A2( _z2[45] ), .A3( n13 ), .Z( _y[45] ) );
XOR3UD1BWP30P140 U77 ( .A1( _z1[46] ), .A2( _z2[46] ), .A3( n14 ), .Z( _y[46] ) );
XOR3UD1BWP30P140 U78 ( .A1( _z1[47] ), .A2( _z2[47] ), .A3( n15 ), .Z( _y[47] ) );
XOR3UD1BWP30P140 U79 ( .A1( _z1[48] ), .A2( _z2[48] ), .A3( n16 ), .Z( _y[48] ) );
XOR3UD1BWP30P140 U80 ( .A1( _z1[49] ), .A2( _z2[49] ), .A3( n17 ), .Z( _y[49] ) );
XOR3UD1BWP30P140 U81 ( .A1( _z1[50] ), .A2( _z2[50] ), .A3( n18 ), .Z( _y[50] ) );
XOR3UD1BWP30P140 U82 ( .A1( _z1[51] ), .A2( _z2[51] ), .A3( n19 ), .Z( _y[51] ) );
XOR3UD1BWP30P140 U83 ( .A1( _z1[52] ), .A2( _z2[52] ), .A3( n20 ), .Z( _y[52] ) );
XOR3UD1BWP30P140 U84 ( .A1( _z1[53] ), .A2( _z2[53] ), .A3( n21 ), .Z( _y[53] ) );
XOR3UD1BWP30P140 U85 ( .A1( _z1[54] ), .A2( _z2[54] ), .A3( n22 ), .Z( _y[54] ) );
XOR3UD1BWP30P140 U86 ( .A1( _z1[55] ), .A2( _z2[55] ), .A3( n23 ), .Z( _y[55] ) );
XOR3UD1BWP30P140 U87 ( .A1( _z1[56] ), .A2( _z2[56] ), .A3( n24 ), .Z( _y[56] ) );
XOR3UD1BWP30P140 U88 ( .A1( _z1[57] ), .A2( _z2[57] ), .A3( n25 ), .Z( _y[57] ) );
XOR3UD1BWP30P140 U89 ( .A1( _z1[58] ), .A2( _z2[58] ), .A3( n26 ), .Z( _y[58] ) );
XOR3UD1BWP30P140 U90 ( .A1( _z1[59] ), .A2( _z2[59] ), .A3( n27 ), .Z( _y[59] ) );
XOR3UD1BWP30P140 U91 ( .A1( _z1[60] ), .A2( _z2[60] ), .A3( n28 ), .Z( _y[60] ) );
XOR3UD1BWP30P140 U92 ( .A1( _z1[61] ), .A2( _z2[61] ), .A3( n29 ), .Z( _y[61] ) );
XOR3UD1BWP30P140 U93 ( .A1( _z1[62] ), .A2( _z2[62] ), .A3( n30 ), .Z( _y[62] ) );
endmodule
