module gf_mul_128_0 ( a, b, C_g1, rst_n, c );
input [127:0] a;
input [127:0] b;
input [21:0] C_g1;
input rst_n;
output [127:0] c;
wire [254:0] d;
assign _a[0] = a[0];
assign _a[1] = a[1];
assign _a[2] = a[2];
assign _a[3] = a[3];
assign _a[4] = a[4];
assign _a[5] = a[5];
assign _a[6] = a[6];
assign _a[7] = a[7];
assign _a[8] = a[8];
assign _a[9] = a[9];
assign _a[10] = a[10];
assign _a[11] = a[11];
assign _a[12] = a[12];
assign _a[13] = a[13];
assign _a[14] = a[14];
assign _a[15] = a[15];
assign _a[16] = a[16];
assign _a[17] = a[17];
assign _a[18] = a[18];
assign _a[19] = a[19];
assign _a[20] = a[20];
assign _a[21] = a[21];
assign _a[22] = a[22];
assign _a[23] = a[23];
assign _a[24] = a[24];
assign _a[25] = a[25];
assign _a[26] = a[26];
assign _a[27] = a[27];
assign _a[28] = a[28];
assign _a[29] = a[29];
assign _a[30] = a[30];
assign _a[31] = a[31];
assign _a[32] = a[32];
assign _a[33] = a[33];
assign _a[34] = a[34];
assign _a[35] = a[35];
assign _a[36] = a[36];
assign _a[37] = a[37];
assign _a[38] = a[38];
assign _a[39] = a[39];
assign _a[40] = a[40];
assign _a[41] = a[41];
assign _a[42] = a[42];
assign _a[43] = a[43];
assign _a[44] = a[44];
assign _a[45] = a[45];
assign _a[46] = a[46];
assign _a[47] = a[47];
assign _a[48] = a[48];
assign _a[49] = a[49];
assign _a[50] = a[50];
assign _a[51] = a[51];
assign _a[52] = a[52];
assign _a[53] = a[53];
assign _a[54] = a[54];
assign _a[55] = a[55];
assign _a[56] = a[56];
assign _a[57] = a[57];
assign _a[58] = a[58];
assign _a[59] = a[59];
assign _a[60] = a[60];
assign _a[61] = a[61];
assign _a[62] = a[62];
assign _a[63] = a[63];
assign _a[64] = a[64];
assign _a[65] = a[65];
assign _a[66] = a[66];
assign _a[67] = a[67];
assign _a[68] = a[68];
assign _a[69] = a[69];
assign _a[70] = a[70];
assign _a[71] = a[71];
assign _a[72] = a[72];
assign _a[73] = a[73];
assign _a[74] = a[74];
assign _a[75] = a[75];
assign _a[76] = a[76];
assign _a[77] = a[77];
assign _a[78] = a[78];
assign _a[79] = a[79];
assign _a[80] = a[80];
assign _a[81] = a[81];
assign _a[82] = a[82];
assign _a[83] = a[83];
assign _a[84] = a[84];
assign _a[85] = a[85];
assign _a[86] = a[86];
assign _a[87] = a[87];
assign _a[88] = a[88];
assign _a[89] = a[89];
assign _a[90] = a[90];
assign _a[91] = a[91];
assign _a[92] = a[92];
assign _a[93] = a[93];
assign _a[94] = a[94];
assign _a[95] = a[95];
assign _a[96] = a[96];
assign _a[97] = a[97];
assign _a[98] = a[98];
assign _a[99] = a[99];
assign _a[100] = a[100];
assign _a[101] = a[101];
assign _a[102] = a[102];
assign _a[103] = a[103];
assign _a[104] = a[104];
assign _a[105] = a[105];
assign _a[106] = a[106];
assign _a[107] = a[107];
assign _a[108] = a[108];
assign _a[109] = a[109];
assign _a[110] = a[110];
assign _a[111] = a[111];
assign _a[112] = a[112];
assign _a[113] = a[113];
assign _a[114] = a[114];
assign _a[115] = a[115];
assign _a[116] = a[116];
assign _a[117] = a[117];
assign _a[118] = a[118];
assign _a[119] = a[119];
assign _a[120] = a[120];
assign _a[121] = a[121];
assign _a[122] = a[122];
assign _a[123] = a[123];
assign _a[124] = a[124];
assign _a[125] = a[125];
assign _a[126] = a[126];
assign _a[127] = a[127];
assign _b[0] = b[0];
assign _b[1] = b[1];
assign _b[2] = b[2];
assign _b[3] = b[3];
assign _b[4] = b[4];
assign _b[5] = b[5];
assign _b[6] = b[6];
assign _b[7] = b[7];
assign _b[8] = b[8];
assign _b[9] = b[9];
assign _b[10] = b[10];
assign _b[11] = b[11];
assign _b[12] = b[12];
assign _b[13] = b[13];
assign _b[14] = b[14];
assign _b[15] = b[15];
assign _b[16] = b[16];
assign _b[17] = b[17];
assign _b[18] = b[18];
assign _b[19] = b[19];
assign _b[20] = b[20];
assign _b[21] = b[21];
assign _b[22] = b[22];
assign _b[23] = b[23];
assign _b[24] = b[24];
assign _b[25] = b[25];
assign _b[26] = b[26];
assign _b[27] = b[27];
assign _b[28] = b[28];
assign _b[29] = b[29];
assign _b[30] = b[30];
assign _b[31] = b[31];
assign _b[32] = b[32];
assign _b[33] = b[33];
assign _b[34] = b[34];
assign _b[35] = b[35];
assign _b[36] = b[36];
assign _b[37] = b[37];
assign _b[38] = b[38];
assign _b[39] = b[39];
assign _b[40] = b[40];
assign _b[41] = b[41];
assign _b[42] = b[42];
assign _b[43] = b[43];
assign _b[44] = b[44];
assign _b[45] = b[45];
assign _b[46] = b[46];
assign _b[47] = b[47];
assign _b[48] = b[48];
assign _b[49] = b[49];
assign _b[50] = b[50];
assign _b[51] = b[51];
assign _b[52] = b[52];
assign _b[53] = b[53];
assign _b[54] = b[54];
assign _b[55] = b[55];
assign _b[56] = b[56];
assign _b[57] = b[57];
assign _b[58] = b[58];
assign _b[59] = b[59];
assign _b[60] = b[60];
assign _b[61] = b[61];
assign _b[62] = b[62];
assign _b[63] = b[63];
assign _b[64] = b[64];
assign _b[65] = b[65];
assign _b[66] = b[66];
assign _b[67] = b[67];
assign _b[68] = b[68];
assign _b[69] = b[69];
assign _b[70] = b[70];
assign _b[71] = b[71];
assign _b[72] = b[72];
assign _b[73] = b[73];
assign _b[74] = b[74];
assign _b[75] = b[75];
assign _b[76] = b[76];
assign _b[77] = b[77];
assign _b[78] = b[78];
assign _b[79] = b[79];
assign _b[80] = b[80];
assign _b[81] = b[81];
assign _b[82] = b[82];
assign _b[83] = b[83];
assign _b[84] = b[84];
assign _b[85] = b[85];
assign _b[86] = b[86];
assign _b[87] = b[87];
assign _b[88] = b[88];
assign _b[89] = b[89];
assign _b[90] = b[90];
assign _b[91] = b[91];
assign _b[92] = b[92];
assign _b[93] = b[93];
assign _b[94] = b[94];
assign _b[95] = b[95];
assign _b[96] = b[96];
assign _b[97] = b[97];
assign _b[98] = b[98];
assign _b[99] = b[99];
assign _b[100] = b[100];
assign _b[101] = b[101];
assign _b[102] = b[102];
assign _b[103] = b[103];
assign _b[104] = b[104];
assign _b[105] = b[105];
assign _b[106] = b[106];
assign _b[107] = b[107];
assign _b[108] = b[108];
assign _b[109] = b[109];
assign _b[110] = b[110];
assign _b[111] = b[111];
assign _b[112] = b[112];
assign _b[113] = b[113];
assign _b[114] = b[114];
assign _b[115] = b[115];
assign _b[116] = b[116];
assign _b[117] = b[117];
assign _b[118] = b[118];
assign _b[119] = b[119];
assign _b[120] = b[120];
assign _b[121] = b[121];
assign _b[122] = b[122];
assign _b[123] = b[123];
assign _b[124] = b[124];
assign _b[125] = b[125];
assign _b[126] = b[126];
assign _b[127] = b[127];
assign _C_g1[0] = C_g1[0];
assign _C_g1[1] = C_g1[1];
assign _C_g1[2] = C_g1[2];
assign _C_g1[3] = C_g1[3];
assign _C_g1[4] = C_g1[4];
assign _C_g1[5] = C_g1[5];
assign _C_g1[6] = C_g1[6];
assign _C_g1[7] = C_g1[7];
assign _C_g1[8] = C_g1[8];
assign _C_g1[9] = C_g1[9];
assign _C_g1[10] = C_g1[10];
assign _C_g1[11] = C_g1[11];
assign _C_g1[12] = C_g1[12];
assign _C_g1[13] = C_g1[13];
assign _C_g1[14] = C_g1[14];
assign _C_g1[15] = C_g1[15];
assign _C_g1[16] = C_g1[16];
assign _C_g1[17] = C_g1[17];
assign _C_g1[18] = C_g1[18];
assign _C_g1[19] = C_g1[19];
assign _C_g1[20] = C_g1[20];
assign _C_g1[21] = C_g1[21];
assign _rst_n = rst_n;
assign c[0] = _c[0];
assign c[1] = _c[1];
assign c[2] = _c[2];
assign c[3] = _c[3];
assign c[4] = _c[4];
assign c[5] = _c[5];
assign c[6] = _c[6];
assign c[7] = _c[7];
assign c[8] = _c[8];
assign c[9] = _c[9];
assign c[10] = _c[10];
assign c[11] = _c[11];
assign c[12] = _c[12];
assign c[13] = _c[13];
assign c[14] = _c[14];
assign c[15] = _c[15];
assign c[16] = _c[16];
assign c[17] = _c[17];
assign c[18] = _c[18];
assign c[19] = _c[19];
assign c[20] = _c[20];
assign c[21] = _c[21];
assign c[22] = _c[22];
assign c[23] = _c[23];
assign c[24] = _c[24];
assign c[25] = _c[25];
assign c[26] = _c[26];
assign c[27] = _c[27];
assign c[28] = _c[28];
assign c[29] = _c[29];
assign c[30] = _c[30];
assign c[31] = _c[31];
assign c[32] = _c[32];
assign c[33] = _c[33];
assign c[34] = _c[34];
assign c[35] = _c[35];
assign c[36] = _c[36];
assign c[37] = _c[37];
assign c[38] = _c[38];
assign c[39] = _c[39];
assign c[40] = _c[40];
assign c[41] = _c[41];
assign c[42] = _c[42];
assign c[43] = _c[43];
assign c[44] = _c[44];
assign c[45] = _c[45];
assign c[46] = _c[46];
assign c[47] = _c[47];
assign c[48] = _c[48];
assign c[49] = _c[49];
assign c[50] = _c[50];
assign c[51] = _c[51];
assign c[52] = _c[52];
assign c[53] = _c[53];
assign c[54] = _c[54];
assign c[55] = _c[55];
assign c[56] = _c[56];
assign c[57] = _c[57];
assign c[58] = _c[58];
assign c[59] = _c[59];
assign c[60] = _c[60];
assign c[61] = _c[61];
assign c[62] = _c[62];
assign c[63] = _c[63];
assign c[64] = _c[64];
assign c[65] = _c[65];
assign c[66] = _c[66];
assign c[67] = _c[67];
assign c[68] = _c[68];
assign c[69] = _c[69];
assign c[70] = _c[70];
assign c[71] = _c[71];
assign c[72] = _c[72];
assign c[73] = _c[73];
assign c[74] = _c[74];
assign c[75] = _c[75];
assign c[76] = _c[76];
assign c[77] = _c[77];
assign c[78] = _c[78];
assign c[79] = _c[79];
assign c[80] = _c[80];
assign c[81] = _c[81];
assign c[82] = _c[82];
assign c[83] = _c[83];
assign c[84] = _c[84];
assign c[85] = _c[85];
assign c[86] = _c[86];
assign c[87] = _c[87];
assign c[88] = _c[88];
assign c[89] = _c[89];
assign c[90] = _c[90];
assign c[91] = _c[91];
assign c[92] = _c[92];
assign c[93] = _c[93];
assign c[94] = _c[94];
assign c[95] = _c[95];
assign c[96] = _c[96];
assign c[97] = _c[97];
assign c[98] = _c[98];
assign c[99] = _c[99];
assign c[100] = _c[100];
assign c[101] = _c[101];
assign c[102] = _c[102];
assign c[103] = _c[103];
assign c[104] = _c[104];
assign c[105] = _c[105];
assign c[106] = _c[106];
assign c[107] = _c[107];
assign c[108] = _c[108];
assign c[109] = _c[109];
assign c[110] = _c[110];
assign c[111] = _c[111];
assign c[112] = _c[112];
assign c[113] = _c[113];
assign c[114] = _c[114];
assign c[115] = _c[115];
assign c[116] = _c[116];
assign c[117] = _c[117];
assign c[118] = _c[118];
assign c[119] = _c[119];
assign c[120] = _c[120];
assign c[121] = _c[121];
assign c[122] = _c[122];
assign c[123] = _c[123];
assign c[124] = _c[124];
assign c[125] = _c[125];
assign c[126] = _c[126];
assign c[127] = _c[127];
OKA_128bit_0 mul_128_x ( .a( _a ), 
.b( _b ), 
.y( d ), 
.C_g1( _C_g1 ), 
.rst_n( _rst_n ) );
reduction_0 reduction_x ( .a( d ), 
.C_g1( _C_g1 ), 
.rst_n( _rst_n ), 
.b( _c ) );
endmodule
