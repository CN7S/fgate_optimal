module XOR2UD1BWP30P140 (
    A1,A2,Z
);
    input A1;
    input A2;
    output Z;
endmodule

module XOR3UD1BWP30P140 (
    A1,A2,A3,Z
);
    input A1;
    input A2;
    input A3;
    output Z;
endmodule
module XOR4D1BWP30P140 (
    A1,A2,A3,A4,Z
);
    input A1;
    input A2;
    input A3;
    input A4;
    output Z;
endmodule

module CKND2D1BWP30P140 (
    A1,A2,ZN
);
    input A1;
    input A2;
    output ZN;
endmodule

module NR2D1BWP30P140 (
    A1,A2,ZN
);
    input A1;
    input A2;
    output ZN;
endmodule
module AN2D1BWP30P140 (
    A1,A2,Z
);
    input A1;
    input A2;
    output Z;
endmodule
module INR2D1BWP30P140 (
    A1,B1,ZN
);
    input A1;
    input B1;
    output ZN;
endmodule
module INVD1BWP30P140 (
    I,ZN
);
    input I;
    output ZN;
endmodule
module XNR3UD1BWP30P140 (
    A1,A2,A3,ZN
);
    input A1,A2,A3;
    output ZN;
endmodule

module XNR2UD1BWP30P140 (
    A1,A2,ZN
);
    input A1,A2;
    output ZN;
endmodule