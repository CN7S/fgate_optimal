module gf_mul_128 ( a, b, c, C_g1, rst_n );
  input [127:0] a;
  input [127:0] b;
  input [21:0] C_g1;
  input rst_n;
  output [127:0] c;

  wire   [254:0] d;


  OKA_128bit mul_128_x ( .a({a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7],
        a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17],
        a[18], a[19], a[20], a[21], a[22], a[23], a[24], a[25], a[26], a[27],
        a[28], a[29], a[30], a[31], a[32], a[33], a[34], a[35], a[36], a[37],
        a[38], a[39], a[40], a[41], a[42], a[43], a[44], a[45], a[46], a[47],
        a[48], a[49], a[50], a[51], a[52], a[53], a[54], a[55], a[56], a[57],
        a[58], a[59], a[60], a[61], a[62], a[63], a[64], a[65], a[66], a[67],
        a[68], a[69], a[70], a[71], a[72], a[73], a[74], a[75], a[76], a[77],
        a[78], a[79], a[80], a[81], a[82], a[83], a[84], a[85], a[86], a[87],
        a[88], a[89], a[90], a[91], a[92], a[93], a[94], a[95], a[96], a[97],
        a[98], a[99], a[100], a[101], a[102], a[103], a[104], a[105], a[106],
        a[107], a[108], a[109], a[110], a[111], a[112], a[113], a[114], a[115],
        a[116], a[117], a[118], a[119], a[120], a[121], a[122], a[123], a[124],
        a[125], a[126], a[127]}), .b({b[0], b[1], b[2], b[3], b[4], b[5], b[6],
        b[7], b[8], b[9], b[10], b[11], b[12], b[13], b[14], b[15], b[16],
        b[17], b[18], b[19], b[20], b[21], b[22], b[23], b[24], b[25], b[26],
        b[27], b[28], b[29], b[30], b[31], b[32], b[33], b[34], b[35], b[36],
        b[37], b[38], b[39], b[40], b[41], b[42], b[43], b[44], b[45], b[46],
        b[47], b[48], b[49], b[50], b[51], b[52], b[53], b[54], b[55], b[56],
        b[57], b[58], b[59], b[60], b[61], b[62], b[63], b[64], b[65], b[66],
        b[67], b[68], b[69], b[70], b[71], b[72], b[73], b[74], b[75], b[76],
        b[77], b[78], b[79], b[80], b[81], b[82], b[83], b[84], b[85], b[86],
        b[87], b[88], b[89], b[90], b[91], b[92], b[93], b[94], b[95], b[96],
        b[97], b[98], b[99], b[100], b[101], b[102], b[103], b[104], b[105],
        b[106], b[107], b[108], b[109], b[110], b[111], b[112], b[113], b[114],
        b[115], b[116], b[117], b[118], b[119], b[120], b[121], b[122], b[123],
        b[124], b[125], b[126], b[127]}), .y(d), .C_g1(C_g1), .rst_n(rst_n) );

  reduction reduction_x ( .a(d), .b({c[0], c[1], c[2], c[3], c[4], c[5],
        c[6], c[7], c[8], c[9], c[10], c[11], c[12], c[13], c[14], c[15],
        c[16], c[17], c[18], c[19], c[20], c[21], c[22], c[23], c[24], c[25],
        c[26], c[27], c[28], c[29], c[30], c[31], c[32], c[33], c[34], c[35],
        c[36], c[37], c[38], c[39], c[40], c[41], c[42], c[43], c[44], c[45],
        c[46], c[47], c[48], c[49], c[50], c[51], c[52], c[53], c[54], c[55],
        c[56], c[57], c[58], c[59], c[60], c[61], c[62], c[63], c[64], c[65],
        c[66], c[67], c[68], c[69], c[70], c[71], c[72], c[73], c[74], c[75],
        c[76], c[77], c[78], c[79], c[80], c[81], c[82], c[83], c[84], c[85],
        c[86], c[87], c[88], c[89], c[90], c[91], c[92], c[93], c[94], c[95],
        c[96], c[97], c[98], c[99], c[100], c[101], c[102], c[103], c[104],
        c[105], c[106], c[107], c[108], c[109], c[110], c[111], c[112], c[113],
        c[114], c[115], c[116], c[117], c[118], c[119], c[120], c[121], c[122],
        c[123], c[124], c[125], c[126], c[127]}),
        .C_g1(C_g1), .rst_n(rst_n) );
endmodule
