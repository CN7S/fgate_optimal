module os_16bit_21 ( z0, z1, z2, o, y );
input [7:0] z0;
input [14:0] z1;
input [7:0] z2;
input [6:0] o;
output [14:0] y;
wire [7:0] _z0;
wire [14:0] _z1;
wire [7:0] _z2;
wire [6:0] _o;
wire [14:0] _y;
assign _z0 = z0;
assign _z1 = z1;
assign _z2 = z2;
assign _o = o;
assign y = _y;
XOR3UD1BWP30P140 U7 ( .A1( _z1[0] ), .A2( _z0[0] ), .A3( _o[0] ), .Z( _y[0] ) );
XOR3UD1BWP30P140 U8 ( .A1( _z1[1] ), .A2( _z0[1] ), .A3( _o[1] ), .Z( _y[1] ) );
XOR3UD1BWP30P140 U9 ( .A1( _z1[2] ), .A2( _z0[2] ), .A3( _o[2] ), .Z( _y[2] ) );
XOR3UD1BWP30P140 U10 ( .A1( _z1[3] ), .A2( _z0[3] ), .A3( _o[3] ), .Z( _y[3] ) );
XOR3UD1BWP30P140 U11 ( .A1( _z1[4] ), .A2( _z0[4] ), .A3( _o[4] ), .Z( _y[4] ) );
XOR3UD1BWP30P140 U12 ( .A1( _z1[5] ), .A2( _z0[5] ), .A3( _o[5] ), .Z( _y[5] ) );
XOR3UD1BWP30P140 U13 ( .A1( _z1[6] ), .A2( _z0[6] ), .A3( _o[6] ), .Z( _y[6] ) );
XOR3UD1BWP30P140 U14 ( .A1( _z2[0] ), .A2( _z1[7] ), .A3( _z0[7] ), .Z( _y[7] ) );
XOR3UD1BWP30P140 U15 ( .A1( _z1[8] ), .A2( _z2[1] ), .A3( _o[0] ), .Z( _y[8] ) );
XOR3UD1BWP30P140 U16 ( .A1( _z1[9] ), .A2( _z2[2] ), .A3( _o[1] ), .Z( _y[9] ) );
XOR3UD1BWP30P140 U17 ( .A1( _z1[10] ), .A2( _z2[3] ), .A3( _o[2] ), .Z( _y[10] ) );
XOR3UD1BWP30P140 U18 ( .A1( _z1[11] ), .A2( _z2[4] ), .A3( _o[3] ), .Z( _y[11] ) );
XOR3UD1BWP30P140 U19 ( .A1( _z1[12] ), .A2( _z2[5] ), .A3( _o[4] ), .Z( _y[12] ) );
XOR3UD1BWP30P140 U20 ( .A1( _z1[13] ), .A2( _z2[6] ), .A3( _o[5] ), .Z( _y[13] ) );
XOR3UD1BWP30P140 U21 ( .A1( _z1[14] ), .A2( _z2[7] ), .A3( _o[6] ), .Z( _y[14] ) );
endmodule
