module reduction ( a, b );
input [254:0] a;
output [127:0] b;
wire [127:0] _b;
wire [254:0] _a;
wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34, n35, n36, n37, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50, n52, n53, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145;
assign _a = a;
assign b = _b;
XOR2UD1BWP30P140 U1 ( .A1( _a[252] ), .A2( _a[131] ), .Z( n97 ) );
XOR2UD1BWP30P140 U2 ( .A1( _a[253] ), .A2( _a[254] ), .Z( n98 ) );
XOR2UD1BWP30P140 U3 ( .A1( _a[132] ), .A2( _a[253] ), .Z( n104 ) );
XOR2UD1BWP30P140 U4 ( .A1( _a[129] ), .A2( _a[250] ), .Z( n76 ) );
XOR2UD1BWP30P140 U5 ( .A1( n6 ), .A2( _a[240] ), .Z( n139 ) );
XNR2UD1BWP30P140 U6 ( .A1( _a[250] ), .A2( _a[251] ), .ZN( n118 ) );
XOR2UD1BWP30P140 U7 ( .A1( n7 ), .A2( _a[238] ), .Z( n140 ) );
XOR2UD1BWP30P140 U8 ( .A1( n8 ), .A2( _a[236] ), .Z( n141 ) );
XOR2UD1BWP30P140 U9 ( .A1( n9 ), .A2( _a[234] ), .Z( n142 ) );
XOR2UD1BWP30P140 U10 ( .A1( n10 ), .A2( _a[232] ), .Z( n143 ) );
XOR2UD1BWP30P140 U11 ( .A1( n11 ), .A2( _a[230] ), .Z( n144 ) );
XOR2UD1BWP30P140 U12 ( .A1( n12 ), .A2( _a[228] ), .Z( n145 ) );
XOR2UD1BWP30P140 U13 ( .A1( n14 ), .A2( _a[226] ), .Z( n69 ) );
XNR2UD1BWP30P140 U14 ( .A1( _a[163] ), .A2( _a[164] ), .ZN( n113 ) );
XOR2UD1BWP30P140 U15 ( .A1( _a[133] ), .A2( _a[134] ), .Z( n82 ) );
XOR2UD1BWP30P140 U16 ( .A1( _a[135] ), .A2( _a[136] ), .Z( n67 ) );
XOR2UD1BWP30P140 U17 ( .A1( _a[139] ), .A2( _a[140] ), .Z( n130 ) );
XNR2UD1BWP30P140 U18 ( .A1( _a[186] ), .A2( _a[187] ), .ZN( n96 ) );
XOR2UD1BWP30P140 U19 ( .A1( n16 ), .A2( _a[224] ), .Z( n71 ) );
XNR2UD1BWP30P140 U20 ( .A1( _a[241] ), .A2( _a[242] ), .ZN( n138 ) );
XOR2UD1BWP30P140 U21 ( .A1( n19 ), .A2( _a[214] ), .Z( n78 ) );
XOR2UD1BWP30P140 U22 ( .A1( n22 ), .A2( _a[208] ), .Z( n81 ) );
XOR2UD1BWP30P140 U23 ( .A1( n29 ), .A2( _a[196] ), .Z( n90 ) );
XOR2UD1BWP30P140 U24 ( .A1( n30 ), .A2( _a[194] ), .Z( n92 ) );
XOR2UD1BWP30P140 U25 ( .A1( n23 ), .A2( _a[206] ), .Z( n84 ) );
XOR2UD1BWP30P140 U26 ( .A1( n24 ), .A2( _a[204] ), .Z( n85 ) );
XOR2UD1BWP30P140 U27 ( .A1( n25 ), .A2( _a[202] ), .Z( n86 ) );
XOR2UD1BWP30P140 U28 ( .A1( n26 ), .A2( _a[200] ), .Z( n87 ) );
XOR2UD1BWP30P140 U29 ( .A1( n27 ), .A2( _a[198] ), .Z( n88 ) );
XOR2UD1BWP30P140 U30 ( .A1( n18 ), .A2( _a[216] ), .Z( n77 ) );
XOR2UD1BWP30P140 U31 ( .A1( n20 ), .A2( _a[212] ), .Z( n79 ) );
XOR2UD1BWP30P140 U32 ( .A1( n21 ), .A2( _a[210] ), .Z( n80 ) );
XNR2UD1BWP30P140 U33 ( .A1( n83 ), .A2( _a[254] ), .ZN( n117 ) );
XOR2UD1BWP30P140 U34 ( .A1( n17 ), .A2( _a[222] ), .Z( n73 ) );
XOR2UD1BWP30P140 U35 ( .A1( n31 ), .A2( _a[192] ), .Z( n93 ) );
XOR2UD1BWP30P140 U36 ( .A1( n43 ), .A2( _a[160] ), .Z( n115 ) );
XOR2UD1BWP30P140 U37 ( .A1( n44 ), .A2( _a[158] ), .Z( n116 ) );
XOR2UD1BWP30P140 U38 ( .A1( n45 ), .A2( _a[156] ), .Z( n119 ) );
XOR2UD1BWP30P140 U39 ( .A1( n46 ), .A2( _a[154] ), .Z( n120 ) );
XOR2UD1BWP30P140 U40 ( .A1( n47 ), .A2( _a[152] ), .Z( n121 ) );
XOR2UD1BWP30P140 U41 ( .A1( n48 ), .A2( _a[150] ), .Z( n122 ) );
XOR2UD1BWP30P140 U42 ( .A1( n50 ), .A2( _a[148] ), .Z( n123 ) );
XOR2UD1BWP30P140 U43 ( .A1( n52 ), .A2( _a[146] ), .Z( n125 ) );
XOR2UD1BWP30P140 U44 ( .A1( n53 ), .A2( _a[144] ), .Z( n127 ) );
XNR2UD1BWP30P140 U45 ( .A1( _a[219] ), .A2( _a[220] ), .ZN( n74 ) );
XNR2UD1BWP30P140 U46 ( .A1( _a[217] ), .A2( _a[218] ), .ZN( n75 ) );
XOR2UD1BWP30P140 U47 ( .A1( _a[130] ), .A2( _a[251] ), .Z( n68 ) );
XNR2UD1BWP30P140 U48 ( .A1( _a[243] ), .A2( _a[244] ), .ZN( n137 ) );
XNR2UD1BWP30P140 U49 ( .A1( _a[161] ), .A2( _a[162] ), .ZN( n114 ) );
XNR2UD1BWP30P140 U50 ( .A1( _a[141] ), .A2( _a[142] ), .ZN( n128 ) );
XNR2UD1BWP30P140 U51 ( .A1( _a[189] ), .A2( _a[190] ), .ZN( n94 ) );
XOR2UD1BWP30P140 U52 ( .A1( n34 ), .A2( _a[181] ), .Z( n101 ) );
XOR2UD1BWP30P140 U53 ( .A1( n37 ), .A2( _a[175] ), .Z( n105 ) );
XOR2UD1BWP30P140 U54 ( .A1( n39 ), .A2( _a[173] ), .Z( n106 ) );
XOR2UD1BWP30P140 U55 ( .A1( n40 ), .A2( _a[171] ), .Z( n108 ) );
XOR2UD1BWP30P140 U56 ( .A1( n41 ), .A2( _a[169] ), .Z( n109 ) );
XOR2UD1BWP30P140 U57 ( .A1( n33 ), .A2( _a[183] ), .Z( n100 ) );
XOR2UD1BWP30P140 U58 ( .A1( n35 ), .A2( _a[179] ), .Z( n102 ) );
XOR2UD1BWP30P140 U59 ( .A1( n36 ), .A2( _a[177] ), .Z( n103 ) );
XNR2UD1BWP30P140 U60 ( .A1( _a[246] ), .A2( _a[247] ), .ZN( n134 ) );
XNR2UD1BWP30P140 U61 ( .A1( n98 ), .A2( _a[132] ), .ZN( n89 ) );
XOR2UD1BWP30P140 U62 ( .A1( _a[137] ), .A2( _a[138] ), .Z( n135 ) );
XNR2UD1BWP30P140 U63 ( .A1( _a[184] ), .A2( _a[185] ), .ZN( n99 ) );
XNR2UD1BWP30P140 U64 ( .A1( _a[166] ), .A2( _a[167] ), .ZN( n110 ) );
XNR2UD1BWP30P140 U65 ( .A1( n1 ), .A2( _a[128] ), .ZN( n83 ) );
XOR2UD1BWP30P140 U66 ( .A1( _a[248] ), .A2( n1 ), .Z( n133 ) );
XNR2UD1BWP30P140 U67 ( .A1( _a[0] ), .A2( n117 ), .ZN( _b[0] ) );
INVD1BWP30P140 U68 ( .I( _a[245] ), .ZN( n3 ) );
INVD1BWP30P140 U69 ( .I( _a[249] ), .ZN( n1 ) );
INVD1BWP30P140 U70 ( .I( _a[239] ), .ZN( n6 ) );
INVD1BWP30P140 U71 ( .I( _a[237] ), .ZN( n7 ) );
INVD1BWP30P140 U72 ( .I( _a[235] ), .ZN( n8 ) );
INVD1BWP30P140 U73 ( .I( _a[233] ), .ZN( n9 ) );
INVD1BWP30P140 U74 ( .I( _a[231] ), .ZN( n10 ) );
INVD1BWP30P140 U75 ( .I( _a[229] ), .ZN( n11 ) );
INVD1BWP30P140 U76 ( .I( n107 ), .ZN( _b[45] ) );
XOR4D1BWP30P140 U77 ( .A1( _a[45] ), .A2( _a[171] ), .A3( _a[166] ), .A4( n106 ), .Z( n107 ) );
INVD1BWP30P140 U78 ( .I( n91 ), .ZN( _b[68] ) );
XOR4D1BWP30P140 U79 ( .A1( _a[68] ), .A2( _a[194] ), .A3( _a[189] ), .A4( n90 ), .Z( n91 ) );
INVD1BWP30P140 U80 ( .I( n70 ), .ZN( _b[98] ) );
XOR4D1BWP30P140 U81 ( .A1( _a[98] ), .A2( _a[224] ), .A3( _a[219] ), .A4( n69 ), .Z( n70 ) );
INVD1BWP30P140 U82 ( .I( n72 ), .ZN( _b[96] ) );
XOR4D1BWP30P140 U83 ( .A1( _a[96] ), .A2( _a[222] ), .A3( _a[217] ), .A4( n71 ), .Z( n72 ) );
INVD1BWP30P140 U84 ( .I( _a[182] ), .ZN( n33 ) );
XOR4D1BWP30P140 U85 ( .A1( _a[252] ), .A2( _a[126] ), .A3( _a[247] ), .A4( n98 ), .Z( _b[126] ) );
XOR4D1BWP30P140 U86 ( .A1( _a[252] ), .A2( _a[124] ), .A3( n3 ), .A4( n118 ), .Z( _b[124] ) );
INVD1BWP30P140 U87 ( .I( _a[176] ), .ZN( n36 ) );
INVD1BWP30P140 U88 ( .I( _a[174] ), .ZN( n37 ) );
INVD1BWP30P140 U89 ( .I( _a[170] ), .ZN( n40 ) );
INVD1BWP30P140 U90 ( .I( _a[168] ), .ZN( n41 ) );
INVD1BWP30P140 U91 ( .I( _a[180] ), .ZN( n34 ) );
INVD1BWP30P140 U92 ( .I( _a[178] ), .ZN( n35 ) );
INVD1BWP30P140 U93 ( .I( _a[227] ), .ZN( n12 ) );
INVD1BWP30P140 U94 ( .I( _a[225] ), .ZN( n14 ) );
INVD1BWP30P140 U95 ( .I( _a[223] ), .ZN( n16 ) );
XOR4D1BWP30P140 U96 ( .A1( n65 ), .A2( _a[142] ), .A3( _a[137] ), .A4( n127 ), .Z( _b[16] ) );
INVD1BWP30P140 U97 ( .I( _a[16] ), .ZN( n65 ) );
XOR4D1BWP30P140 U98 ( .A1( n66 ), .A2( n97 ), .A3( _a[133] ), .A4( n89 ), .Z( _b[5] ) );
INVD1BWP30P140 U99 ( .I( _a[5] ), .ZN( n66 ) );
XOR4D1BWP30P140 U100 ( .A1( n63 ), .A2( _a[163] ), .A3( _a[156] ), .A4( n114 ), .Z( _b[35] ) );
INVD1BWP30P140 U101 ( .I( _a[35] ), .ZN( n63 ) );
XOR4D1BWP30P140 U102 ( .A1( n59 ), .A2( _a[186] ), .A3( _a[179] ), .A4( n99 ), .Z( _b[58] ) );
INVD1BWP30P140 U103 ( .I( _a[58] ), .ZN( n59 ) );
XOR4D1BWP30P140 U104 ( .A1( n60 ), .A2( _a[184] ), .A3( _a[177] ), .A4( n100 ), .Z( _b[56] ) );
INVD1BWP30P140 U105 ( .I( _a[56] ), .ZN( n60 ) );
XOR4D1BWP30P140 U106 ( .A1( n64 ), .A2( _a[161] ), .A3( _a[154] ), .A4( n115 ), .Z( _b[33] ) );
INVD1BWP30P140 U107 ( .I( _a[33] ), .ZN( n64 ) );
XOR4D1BWP30P140 U108 ( .A1( n61 ), .A2( _a[169] ), .A3( _a[164] ), .A4( n108 ), .Z( _b[43] ) );
INVD1BWP30P140 U109 ( .I( _a[43] ), .ZN( n61 ) );
XOR4D1BWP30P140 U110 ( .A1( n62 ), .A2( _a[167] ), .A3( _a[162] ), .A4( n109 ), .Z( _b[41] ) );
INVD1BWP30P140 U111 ( .I( _a[41] ), .ZN( n62 ) );
XOR4D1BWP30P140 U112 ( .A1( n58 ), .A2( _a[190] ), .A3( _a[185] ), .A4( n93 ), .Z( _b[64] ) );
INVD1BWP30P140 U113 ( .I( _a[64] ), .ZN( n58 ) );
XOR4D1BWP30P140 U114 ( .A1( n55 ), .A2( _a[219] ), .A3( _a[212] ), .A4( n75 ), .Z( _b[91] ) );
INVD1BWP30P140 U115 ( .I( _a[91] ), .ZN( n55 ) );
XOR4D1BWP30P140 U116 ( .A1( n56 ), .A2( _a[217] ), .A3( _a[210] ), .A4( n77 ), .Z( _b[89] ) );
INVD1BWP30P140 U117 ( .I( _a[89] ), .ZN( n56 ) );
XOR4D1BWP30P140 U118 ( .A1( n2 ), .A2( _a[121] ), .A3( _a[242] ), .A4( n133 ), .Z( _b[121] ) );
INVD1BWP30P140 U119 ( .I( _a[247] ), .ZN( n2 ) );
XOR4D1BWP30P140 U120 ( .A1( n57 ), .A2( _a[192] ), .A3( _a[187] ), .A4( n92 ), .Z( _b[66] ) );
INVD1BWP30P140 U121 ( .I( _a[66] ), .ZN( n57 ) );
XOR4D1BWP30P140 U122 ( .A1( n4 ), .A2( _a[115] ), .A3( _a[236] ), .A4( n138 ), .Z( _b[115] ) );
XOR4D1BWP30P140 U123 ( .A1( n5 ), .A2( _a[113] ), .A3( _a[234] ), .A4( n139 ), .Z( _b[113] ) );
XOR4D1BWP30P140 U124 ( .A1( n7 ), .A2( _a[109] ), .A3( _a[230] ), .A4( n141 ), .Z( _b[109] ) );
XOR4D1BWP30P140 U125 ( .A1( n8 ), .A2( _a[107] ), .A3( _a[228] ), .A4( n142 ), .Z( _b[107] ) );
XOR4D1BWP30P140 U126 ( .A1( n9 ), .A2( _a[105] ), .A3( _a[226] ), .A4( n143 ), .Z( _b[105] ) );
XOR4D1BWP30P140 U127 ( .A1( n10 ), .A2( _a[103] ), .A3( _a[224] ), .A4( n144 ), .Z( _b[103] ) );
XOR4D1BWP30P140 U128 ( .A1( n11 ), .A2( _a[101] ), .A3( _a[222] ), .A4( n145 ), .Z( _b[101] ) );
XOR4D1BWP30P140 U129 ( .A1( n6 ), .A2( _a[111] ), .A3( _a[232] ), .A4( n140 ), .Z( _b[111] ) );
XOR4D1BWP30P140 U130 ( .A1( n1 ), .A2( _a[123] ), .A3( _a[244] ), .A4( n118 ), .Z( _b[123] ) );
XOR4D1BWP30P140 U131 ( .A1( n3 ), .A2( _a[119] ), .A3( _a[240] ), .A4( n134 ), .Z( _b[119] ) );
XOR4D1BWP30P140 U132 ( .A1( n3 ), .A2( _a[117] ), .A3( _a[238] ), .A4( n137 ), .Z( _b[117] ) );
XOR4D1BWP30P140 U133 ( .A1( n136 ), .A2( _a[118] ), .A3( _a[244] ), .A4( _a[239] ), .Z( _b[118] ) );
XNR2UD1BWP30P140 U134 ( .A1( _a[246] ), .A2( n3 ), .ZN( n136 ) );
XOR4D1BWP30P140 U135 ( .A1( _a[250] ), .A2( _a[122] ), .A3( n4 ), .A4( n133 ), .Z( _b[122] ) );
XOR4D1BWP30P140 U136 ( .A1( n112 ), .A2( _a[38] ), .A3( _a[166] ), .A4( _a[165] ), .Z( _b[38] ) );
XOR2UD1BWP30P140 U137 ( .A1( _a[164] ), .A2( _a[159] ), .Z( n112 ) );
XOR4D1BWP30P140 U138 ( .A1( _a[99] ), .A2( n12 ), .A3( _a[220] ), .A4( n69 ), .Z( _b[99] ) );
XOR4D1BWP30P140 U139 ( .A1( _a[97] ), .A2( n14 ), .A3( _a[218] ), .A4( n71 ), .Z( _b[97] ) );
XOR4D1BWP30P140 U140 ( .A1( _a[93] ), .A2( n17 ), .A3( _a[214] ), .A4( n74 ), .Z( _b[93] ) );
XOR4D1BWP30P140 U141 ( .A1( _a[73] ), .A2( n25 ), .A3( _a[194] ), .A4( n87 ), .Z( _b[73] ) );
XOR4D1BWP30P140 U142 ( .A1( _a[69] ), .A2( n27 ), .A3( _a[190] ), .A4( n90 ), .Z( _b[69] ) );
XOR4D1BWP30P140 U143 ( .A1( _a[67] ), .A2( _a[195] ), .A3( n32 ), .A4( n92 ), .Z( _b[67] ) );
XOR4D1BWP30P140 U144 ( .A1( _a[65] ), .A2( n30 ), .A3( _a[186] ), .A4( n93 ), .Z( _b[65] ) );
XOR4D1BWP30P140 U145 ( .A1( _a[95] ), .A2( n16 ), .A3( _a[216] ), .A4( n73 ), .Z( _b[95] ) );
XOR4D1BWP30P140 U146 ( .A1( _a[87] ), .A2( n18 ), .A3( _a[208] ), .A4( n78 ), .Z( _b[87] ) );
XOR4D1BWP30P140 U147 ( .A1( _a[85] ), .A2( n19 ), .A3( _a[206] ), .A4( n79 ), .Z( _b[85] ) );
XOR4D1BWP30P140 U148 ( .A1( _a[83] ), .A2( n20 ), .A3( _a[204] ), .A4( n80 ), .Z( _b[83] ) );
XOR4D1BWP30P140 U149 ( .A1( _a[81] ), .A2( n21 ), .A3( _a[202] ), .A4( n81 ), .Z( _b[81] ) );
XOR4D1BWP30P140 U150 ( .A1( _a[79] ), .A2( n22 ), .A3( _a[200] ), .A4( n84 ), .Z( _b[79] ) );
XOR4D1BWP30P140 U151 ( .A1( _a[77] ), .A2( n23 ), .A3( _a[198] ), .A4( n85 ), .Z( _b[77] ) );
XOR4D1BWP30P140 U152 ( .A1( _a[75] ), .A2( n24 ), .A3( _a[196] ), .A4( n86 ), .Z( _b[75] ) );
XOR4D1BWP30P140 U153 ( .A1( _a[71] ), .A2( n26 ), .A3( _a[192] ), .A4( n88 ), .Z( _b[71] ) );
XOR4D1BWP30P140 U154 ( .A1( n95 ), .A2( _a[61] ), .A3( _a[189] ), .A4( _a[188] ), .Z( _b[61] ) );
XOR2UD1BWP30P140 U155 ( .A1( _a[187] ), .A2( _a[182] ), .Z( n95 ) );
XOR4D1BWP30P140 U156 ( .A1( _a[63] ), .A2( n31 ), .A3( _a[184] ), .A4( n94 ), .Z( _b[63] ) );
XOR4D1BWP30P140 U157 ( .A1( _a[59] ), .A2( _a[185] ), .A3( n34 ), .A4( n96 ), .Z( _b[59] ) );
XOR4D1BWP30P140 U158 ( .A1( _a[57] ), .A2( _a[183] ), .A3( n35 ), .A4( n99 ), .Z( _b[57] ) );
XOR4D1BWP30P140 U159 ( .A1( _a[55] ), .A2( _a[181] ), .A3( n36 ), .A4( n100 ), .Z( _b[55] ) );
XOR4D1BWP30P140 U160 ( .A1( _a[53] ), .A2( _a[179] ), .A3( n37 ), .A4( n101 ), .Z( _b[53] ) );
XOR4D1BWP30P140 U161 ( .A1( _a[37] ), .A2( n42 ), .A3( _a[158] ), .A4( n113 ), .Z( _b[37] ) );
XOR4D1BWP30P140 U162 ( .A1( _a[51] ), .A2( _a[177] ), .A3( n39 ), .A4( n102 ), .Z( _b[51] ) );
XOR4D1BWP30P140 U163 ( .A1( _a[49] ), .A2( _a[175] ), .A3( n40 ), .A4( n103 ), .Z( _b[49] ) );
XOR4D1BWP30P140 U164 ( .A1( _a[47] ), .A2( _a[173] ), .A3( n41 ), .A4( n105 ), .Z( _b[47] ) );
XOR4D1BWP30P140 U165 ( .A1( _a[39] ), .A2( n42 ), .A3( _a[160] ), .A4( n110 ), .Z( _b[39] ) );
INVD1BWP30P140 U166 ( .I( _a[159] ), .ZN( n43 ) );
XOR4D1BWP30P140 U167 ( .A1( _a[31] ), .A2( n43 ), .A3( _a[152] ), .A4( n116 ), .Z( _b[31] ) );
XOR4D1BWP30P140 U168 ( .A1( _a[29] ), .A2( n44 ), .A3( _a[150] ), .A4( n119 ), .Z( _b[29] ) );
XOR4D1BWP30P140 U169 ( .A1( _a[27] ), .A2( n45 ), .A3( _a[148] ), .A4( n120 ), .Z( _b[27] ) );
XOR4D1BWP30P140 U170 ( .A1( _a[25] ), .A2( n46 ), .A3( _a[146] ), .A4( n121 ), .Z( _b[25] ) );
XOR4D1BWP30P140 U171 ( .A1( _a[23] ), .A2( n47 ), .A3( _a[144] ), .A4( n122 ), .Z( _b[23] ) );
XOR4D1BWP30P140 U172 ( .A1( _a[21] ), .A2( n48 ), .A3( _a[142] ), .A4( n123 ), .Z( _b[21] ) );
XOR4D1BWP30P140 U173 ( .A1( _a[19] ), .A2( n50 ), .A3( _a[140] ), .A4( n125 ), .Z( _b[19] ) );
XOR4D1BWP30P140 U174 ( .A1( _a[17] ), .A2( n52 ), .A3( _a[138] ), .A4( n127 ), .Z( _b[17] ) );
XOR4D1BWP30P140 U175 ( .A1( _a[74] ), .A2( _a[200] ), .A3( n29 ), .A4( n86 ), .Z( _b[74] ) );
XOR4D1BWP30P140 U176 ( .A1( _a[72] ), .A2( _a[198] ), .A3( n30 ), .A4( n87 ), .Z( _b[72] ) );
XOR4D1BWP30P140 U177 ( .A1( _a[94] ), .A2( _a[220] ), .A3( n18 ), .A4( n73 ), .Z( _b[94] ) );
XOR4D1BWP30P140 U178 ( .A1( _a[92] ), .A2( _a[218] ), .A3( n19 ), .A4( n74 ), .Z( _b[92] ) );
XOR4D1BWP30P140 U179 ( .A1( _a[90] ), .A2( _a[216] ), .A3( n20 ), .A4( n75 ), .Z( _b[90] ) );
XOR4D1BWP30P140 U180 ( .A1( _a[88] ), .A2( _a[214] ), .A3( n21 ), .A4( n77 ), .Z( _b[88] ) );
XOR4D1BWP30P140 U181 ( .A1( _a[86] ), .A2( _a[212] ), .A3( n22 ), .A4( n78 ), .Z( _b[86] ) );
XOR4D1BWP30P140 U182 ( .A1( _a[84] ), .A2( _a[210] ), .A3( n23 ), .A4( n79 ), .Z( _b[84] ) );
XOR4D1BWP30P140 U183 ( .A1( _a[82] ), .A2( _a[208] ), .A3( n24 ), .A4( n80 ), .Z( _b[82] ) );
XOR4D1BWP30P140 U184 ( .A1( _a[80] ), .A2( _a[206] ), .A3( n25 ), .A4( n81 ), .Z( _b[80] ) );
XOR4D1BWP30P140 U185 ( .A1( _a[78] ), .A2( _a[204] ), .A3( n26 ), .A4( n84 ), .Z( _b[78] ) );
XOR4D1BWP30P140 U186 ( .A1( _a[76] ), .A2( _a[202] ), .A3( n27 ), .A4( n85 ), .Z( _b[76] ) );
XOR4D1BWP30P140 U187 ( .A1( _a[70] ), .A2( _a[196] ), .A3( n31 ), .A4( n88 ), .Z( _b[70] ) );
XOR4D1BWP30P140 U188 ( .A1( n67 ), .A2( n68 ), .A3( _a[9] ), .A4( _a[137] ), .Z( _b[9] ) );
XOR4D1BWP30P140 U189 ( .A1( n67 ), .A2( n76 ), .A3( _a[8] ), .A4( _a[134] ), .Z( _b[8] ) );
XOR4D1BWP30P140 U190 ( .A1( _a[62] ), .A2( n32 ), .A3( _a[183] ), .A4( n94 ), .Z( _b[62] ) );
XOR4D1BWP30P140 U191 ( .A1( _a[60] ), .A2( n32 ), .A3( _a[181] ), .A4( n96 ), .Z( _b[60] ) );
XOR4D1BWP30P140 U192 ( .A1( _a[54] ), .A2( n33 ), .A3( _a[175] ), .A4( n101 ), .Z( _b[54] ) );
XOR4D1BWP30P140 U193 ( .A1( _a[42] ), .A2( n40 ), .A3( _a[163] ), .A4( n109 ), .Z( _b[42] ) );
XOR4D1BWP30P140 U194 ( .A1( _a[40] ), .A2( n41 ), .A3( _a[161] ), .A4( n110 ), .Z( _b[40] ) );
XOR4D1BWP30P140 U195 ( .A1( n82 ), .A2( n83 ), .A3( _a[7] ), .A4( _a[135] ), .Z( _b[7] ) );
XOR4D1BWP30P140 U196 ( .A1( _a[36] ), .A2( _a[162] ), .A3( n44 ), .A4( n113 ), .Z( _b[36] ) );
XOR4D1BWP30P140 U197 ( .A1( _a[34] ), .A2( _a[160] ), .A3( n45 ), .A4( n114 ), .Z( _b[34] ) );
XOR4D1BWP30P140 U198 ( .A1( _a[52] ), .A2( n34 ), .A3( _a[173] ), .A4( n102 ), .Z( _b[52] ) );
XOR4D1BWP30P140 U199 ( .A1( _a[50] ), .A2( n35 ), .A3( _a[171] ), .A4( n103 ), .Z( _b[50] ) );
XOR4D1BWP30P140 U200 ( .A1( _a[48] ), .A2( n36 ), .A3( _a[169] ), .A4( n105 ), .Z( _b[48] ) );
XOR4D1BWP30P140 U201 ( .A1( _a[46] ), .A2( n37 ), .A3( _a[167] ), .A4( n106 ), .Z( _b[46] ) );
XOR4D1BWP30P140 U202 ( .A1( _a[15] ), .A2( n53 ), .A3( _a[136] ), .A4( n128 ), .Z( _b[15] ) );
XOR4D1BWP30P140 U203 ( .A1( _a[44] ), .A2( _a[172] ), .A3( n42 ), .A4( n108 ), .Z( _b[44] ) );
XOR4D1BWP30P140 U204 ( .A1( n104 ), .A2( n135 ), .A3( _a[139] ), .A4( _a[11] ), .Z( _b[11] ) );
XOR4D1BWP30P140 U205 ( .A1( _a[32] ), .A2( _a[158] ), .A3( n46 ), .A4( n115 ), .Z( _b[32] ) );
XOR4D1BWP30P140 U206 ( .A1( _a[30] ), .A2( _a[156] ), .A3( n47 ), .A4( n116 ), .Z( _b[30] ) );
XOR4D1BWP30P140 U207 ( .A1( _a[28] ), .A2( _a[154] ), .A3( n48 ), .A4( n119 ), .Z( _b[28] ) );
XOR4D1BWP30P140 U208 ( .A1( _a[26] ), .A2( _a[152] ), .A3( n50 ), .A4( n120 ), .Z( _b[26] ) );
XOR4D1BWP30P140 U209 ( .A1( _a[24] ), .A2( _a[150] ), .A3( n52 ), .A4( n121 ), .Z( _b[24] ) );
XOR4D1BWP30P140 U210 ( .A1( _a[22] ), .A2( _a[148] ), .A3( n53 ), .A4( n122 ), .Z( _b[22] ) );
XOR4D1BWP30P140 U211 ( .A1( n132 ), .A2( _a[125] ), .A3( _a[251] ), .A4( _a[246] ), .Z( _b[125] ) );
XOR2UD1BWP30P140 U212 ( .A1( _a[253] ), .A2( _a[252] ), .Z( n132 ) );
XOR4D1BWP30P140 U213 ( .A1( n97 ), .A2( n135 ), .A3( _a[136] ), .A4( _a[10] ), .Z( _b[10] ) );
XOR4D1BWP30P140 U214 ( .A1( n97 ), .A2( n104 ), .A3( _a[4] ), .A4( n68 ), .Z( _b[4] ) );
XOR4D1BWP30P140 U215 ( .A1( _a[242] ), .A2( _a[116] ), .A3( n7 ), .A4( n137 ), .Z( _b[116] ) );
XOR4D1BWP30P140 U216 ( .A1( _a[141] ), .A2( _a[13] ), .A3( _a[134] ), .A4( n130 ), .Z( _b[13] ) );
XOR4D1BWP30P140 U217 ( .A1( _a[238] ), .A2( _a[112] ), .A3( n9 ), .A4( n139 ), .Z( _b[112] ) );
XOR4D1BWP30P140 U218 ( .A1( _a[236] ), .A2( _a[110] ), .A3( n10 ), .A4( n140 ), .Z( _b[110] ) );
XOR4D1BWP30P140 U219 ( .A1( _a[234] ), .A2( _a[108] ), .A3( n11 ), .A4( n141 ), .Z( _b[108] ) );
XOR4D1BWP30P140 U220 ( .A1( _a[232] ), .A2( _a[106] ), .A3( n12 ), .A4( n142 ), .Z( _b[106] ) );
XOR4D1BWP30P140 U221 ( .A1( _a[230] ), .A2( _a[104] ), .A3( n14 ), .A4( n143 ), .Z( _b[104] ) );
XOR4D1BWP30P140 U222 ( .A1( _a[228] ), .A2( _a[102] ), .A3( n16 ), .A4( n144 ), .Z( _b[102] ) );
XOR4D1BWP30P140 U223 ( .A1( _a[226] ), .A2( _a[100] ), .A3( n17 ), .A4( n145 ), .Z( _b[100] ) );
XOR4D1BWP30P140 U224 ( .A1( _a[248] ), .A2( _a[120] ), .A3( n5 ), .A4( n134 ), .Z( _b[120] ) );
XOR4D1BWP30P140 U225 ( .A1( _a[240] ), .A2( _a[114] ), .A3( n8 ), .A4( n138 ), .Z( _b[114] ) );
INVD1BWP30P140 U226 ( .I( _a[172] ), .ZN( n39 ) );
INVD1BWP30P140 U227 ( .I( _a[213] ), .ZN( n19 ) );
INVD1BWP30P140 U228 ( .I( _a[207] ), .ZN( n22 ) );
INVD1BWP30P140 U229 ( .I( _a[193] ), .ZN( n30 ) );
INVD1BWP30P140 U230 ( .I( _a[205] ), .ZN( n23 ) );
INVD1BWP30P140 U231 ( .I( _a[203] ), .ZN( n24 ) );
INVD1BWP30P140 U232 ( .I( _a[201] ), .ZN( n25 ) );
INVD1BWP30P140 U233 ( .I( _a[199] ), .ZN( n26 ) );
INVD1BWP30P140 U234 ( .I( _a[197] ), .ZN( n27 ) );
INVD1BWP30P140 U235 ( .I( _a[215] ), .ZN( n18 ) );
INVD1BWP30P140 U236 ( .I( _a[211] ), .ZN( n20 ) );
INVD1BWP30P140 U237 ( .I( _a[209] ), .ZN( n21 ) );
INVD1BWP30P140 U238 ( .I( _a[221] ), .ZN( n17 ) );
INVD1BWP30P140 U239 ( .I( _a[191] ), .ZN( n31 ) );
INVD1BWP30P140 U240 ( .I( _a[188] ), .ZN( n32 ) );
INVD1BWP30P140 U241 ( .I( _a[243] ), .ZN( n4 ) );
INVD1BWP30P140 U242 ( .I( _a[241] ), .ZN( n5 ) );
INVD1BWP30P140 U243 ( .I( _a[155] ), .ZN( n45 ) );
INVD1BWP30P140 U244 ( .I( _a[153] ), .ZN( n46 ) );
INVD1BWP30P140 U245 ( .I( _a[149] ), .ZN( n48 ) );
INVD1BWP30P140 U246 ( .I( _a[143] ), .ZN( n53 ) );
INVD1BWP30P140 U247 ( .I( _a[157] ), .ZN( n44 ) );
INVD1BWP30P140 U248 ( .I( _a[151] ), .ZN( n47 ) );
INVD1BWP30P140 U249 ( .I( _a[147] ), .ZN( n50 ) );
INVD1BWP30P140 U250 ( .I( _a[145] ), .ZN( n52 ) );
INVD1BWP30P140 U251 ( .I( _a[195] ), .ZN( n29 ) );
INVD1BWP30P140 U252 ( .I( _a[165] ), .ZN( n42 ) );
XNR3UD1BWP30P140 U253 ( .A1( _a[130] ), .A2( _a[129] ), .A3( n118 ), .ZN( n111 ) );
XOR3UD1BWP30P140 U254 ( .A1( _a[248] ), .A2( _a[127] ), .A3( n98 ), .Z( _b[127] ) );
XNR3UD1BWP30P140 U255 ( .A1( _a[2] ), .A2( n111 ), .A3( n117 ), .ZN( _b[2] ) );
XNR3UD1BWP30P140 U256 ( .A1( _a[1] ), .A2( n76 ), .A3( n117 ), .ZN( _b[1] ) );
XNR3UD1BWP30P140 U257 ( .A1( _a[6] ), .A2( n82 ), .A3( n89 ), .ZN( _b[6] ) );
XOR3UD1BWP30P140 U258 ( .A1( _a[3] ), .A2( n97 ), .A3( n111 ), .Z( _b[3] ) );
XOR3UD1BWP30P140 U259 ( .A1( _a[12] ), .A2( n130 ), .A3( n131 ), .Z( _b[12] ) );
XOR3UD1BWP30P140 U260 ( .A1( _a[254] ), .A2( _a[138] ), .A3( _a[133] ), .Z( n131 ) );
INVD1BWP30P140 U261 ( .I( n129 ), .ZN( _b[14] ) );
XOR4D1BWP30P140 U262 ( .A1( _a[14] ), .A2( _a[140] ), .A3( _a[135] ), .A4( n128 ), .Z( n129 ) );
INVD1BWP30P140 U263 ( .I( n124 ), .ZN( _b[20] ) );
XOR4D1BWP30P140 U264 ( .A1( _a[20] ), .A2( _a[146] ), .A3( _a[141] ), .A4( n123 ), .Z( n124 ) );
INVD1BWP30P140 U265 ( .I( n126 ), .ZN( _b[18] ) );
XOR4D1BWP30P140 U266 ( .A1( _a[18] ), .A2( _a[144] ), .A3( _a[139] ), .A4( n125 ), .Z( n126 ) );
endmodule
