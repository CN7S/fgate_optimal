module DEL025D1BWP30P140 (I, Z);
    input I;
    output Z;
endmodule
