module s_128bit ( a, b, aa, bb );
input [127:0] a;
input [127:0] b;
output [63:0] aa;
output [63:0] bb;
wire [127:0] _a;
wire [127:0] _b;
wire [63:0] _aa;
wire [63:0] _bb;
assign _a = a;
assign _b = b;
assign aa = _aa;
assign bb = _bb;
XOR2UD1BWP30P140 U0 ( .A1( _a[0] ), .A2( _a[1] ), .Z( _aa[0] ) );
XOR2UD1BWP30P140 U1 ( .A1( _a[2] ), .A2( _a[3] ), .Z( _aa[1] ) );
XOR2UD1BWP30P140 U2 ( .A1( _a[4] ), .A2( _a[5] ), .Z( _aa[2] ) );
XOR2UD1BWP30P140 U3 ( .A1( _a[6] ), .A2( _a[7] ), .Z( _aa[3] ) );
XOR2UD1BWP30P140 U4 ( .A1( _a[8] ), .A2( _a[9] ), .Z( _aa[4] ) );
XOR2UD1BWP30P140 U5 ( .A1( _a[10] ), .A2( _a[11] ), .Z( _aa[5] ) );
XOR2UD1BWP30P140 U6 ( .A1( _a[12] ), .A2( _a[13] ), .Z( _aa[6] ) );
XOR2UD1BWP30P140 U7 ( .A1( _a[14] ), .A2( _a[15] ), .Z( _aa[7] ) );
XOR2UD1BWP30P140 U8 ( .A1( _a[16] ), .A2( _a[17] ), .Z( _aa[8] ) );
XOR2UD1BWP30P140 U9 ( .A1( _a[18] ), .A2( _a[19] ), .Z( _aa[9] ) );
XOR2UD1BWP30P140 U10 ( .A1( _a[20] ), .A2( _a[21] ), .Z( _aa[10] ) );
XOR2UD1BWP30P140 U11 ( .A1( _a[22] ), .A2( _a[23] ), .Z( _aa[11] ) );
XOR2UD1BWP30P140 U12 ( .A1( _a[24] ), .A2( _a[25] ), .Z( _aa[12] ) );
XOR2UD1BWP30P140 U13 ( .A1( _a[26] ), .A2( _a[27] ), .Z( _aa[13] ) );
XOR2UD1BWP30P140 U14 ( .A1( _a[28] ), .A2( _a[29] ), .Z( _aa[14] ) );
XOR2UD1BWP30P140 U15 ( .A1( _a[30] ), .A2( _a[31] ), .Z( _aa[15] ) );
XOR2UD1BWP30P140 U16 ( .A1( _a[32] ), .A2( _a[33] ), .Z( _aa[16] ) );
XOR2UD1BWP30P140 U17 ( .A1( _a[34] ), .A2( _a[35] ), .Z( _aa[17] ) );
XOR2UD1BWP30P140 U18 ( .A1( _a[36] ), .A2( _a[37] ), .Z( _aa[18] ) );
XOR2UD1BWP30P140 U19 ( .A1( _a[38] ), .A2( _a[39] ), .Z( _aa[19] ) );
XOR2UD1BWP30P140 U20 ( .A1( _a[40] ), .A2( _a[41] ), .Z( _aa[20] ) );
XOR2UD1BWP30P140 U21 ( .A1( _a[42] ), .A2( _a[43] ), .Z( _aa[21] ) );
XOR2UD1BWP30P140 U22 ( .A1( _a[44] ), .A2( _a[45] ), .Z( _aa[22] ) );
XOR2UD1BWP30P140 U23 ( .A1( _a[46] ), .A2( _a[47] ), .Z( _aa[23] ) );
XOR2UD1BWP30P140 U24 ( .A1( _a[48] ), .A2( _a[49] ), .Z( _aa[24] ) );
XOR2UD1BWP30P140 U25 ( .A1( _a[50] ), .A2( _a[51] ), .Z( _aa[25] ) );
XOR2UD1BWP30P140 U26 ( .A1( _a[52] ), .A2( _a[53] ), .Z( _aa[26] ) );
XOR2UD1BWP30P140 U27 ( .A1( _a[54] ), .A2( _a[55] ), .Z( _aa[27] ) );
XOR2UD1BWP30P140 U28 ( .A1( _a[56] ), .A2( _a[57] ), .Z( _aa[28] ) );
XOR2UD1BWP30P140 U29 ( .A1( _a[58] ), .A2( _a[59] ), .Z( _aa[29] ) );
XOR2UD1BWP30P140 U30 ( .A1( _a[60] ), .A2( _a[61] ), .Z( _aa[30] ) );
XOR2UD1BWP30P140 U31 ( .A1( _a[62] ), .A2( _a[63] ), .Z( _aa[31] ) );
XOR2UD1BWP30P140 U32 ( .A1( _a[64] ), .A2( _a[65] ), .Z( _aa[32] ) );
XOR2UD1BWP30P140 U33 ( .A1( _a[66] ), .A2( _a[67] ), .Z( _aa[33] ) );
XOR2UD1BWP30P140 U34 ( .A1( _a[68] ), .A2( _a[69] ), .Z( _aa[34] ) );
XOR2UD1BWP30P140 U35 ( .A1( _a[70] ), .A2( _a[71] ), .Z( _aa[35] ) );
XOR2UD1BWP30P140 U36 ( .A1( _a[72] ), .A2( _a[73] ), .Z( _aa[36] ) );
XOR2UD1BWP30P140 U37 ( .A1( _a[74] ), .A2( _a[75] ), .Z( _aa[37] ) );
XOR2UD1BWP30P140 U38 ( .A1( _a[76] ), .A2( _a[77] ), .Z( _aa[38] ) );
XOR2UD1BWP30P140 U39 ( .A1( _a[78] ), .A2( _a[79] ), .Z( _aa[39] ) );
XOR2UD1BWP30P140 U40 ( .A1( _a[80] ), .A2( _a[81] ), .Z( _aa[40] ) );
XOR2UD1BWP30P140 U41 ( .A1( _a[82] ), .A2( _a[83] ), .Z( _aa[41] ) );
XOR2UD1BWP30P140 U42 ( .A1( _a[84] ), .A2( _a[85] ), .Z( _aa[42] ) );
XOR2UD1BWP30P140 U43 ( .A1( _a[86] ), .A2( _a[87] ), .Z( _aa[43] ) );
XOR2UD1BWP30P140 U44 ( .A1( _a[88] ), .A2( _a[89] ), .Z( _aa[44] ) );
XOR2UD1BWP30P140 U45 ( .A1( _a[90] ), .A2( _a[91] ), .Z( _aa[45] ) );
XOR2UD1BWP30P140 U46 ( .A1( _a[92] ), .A2( _a[93] ), .Z( _aa[46] ) );
XOR2UD1BWP30P140 U47 ( .A1( _a[94] ), .A2( _a[95] ), .Z( _aa[47] ) );
XOR2UD1BWP30P140 U48 ( .A1( _a[96] ), .A2( _a[97] ), .Z( _aa[48] ) );
XOR2UD1BWP30P140 U49 ( .A1( _a[98] ), .A2( _a[99] ), .Z( _aa[49] ) );
XOR2UD1BWP30P140 U50 ( .A1( _a[100] ), .A2( _a[101] ), .Z( _aa[50] ) );
XOR2UD1BWP30P140 U51 ( .A1( _a[102] ), .A2( _a[103] ), .Z( _aa[51] ) );
XOR2UD1BWP30P140 U52 ( .A1( _a[104] ), .A2( _a[105] ), .Z( _aa[52] ) );
XOR2UD1BWP30P140 U53 ( .A1( _a[106] ), .A2( _a[107] ), .Z( _aa[53] ) );
XOR2UD1BWP30P140 U54 ( .A1( _a[108] ), .A2( _a[109] ), .Z( _aa[54] ) );
XOR2UD1BWP30P140 U55 ( .A1( _a[110] ), .A2( _a[111] ), .Z( _aa[55] ) );
XOR2UD1BWP30P140 U56 ( .A1( _a[112] ), .A2( _a[113] ), .Z( _aa[56] ) );
XOR2UD1BWP30P140 U57 ( .A1( _a[114] ), .A2( _a[115] ), .Z( _aa[57] ) );
XOR2UD1BWP30P140 U58 ( .A1( _a[116] ), .A2( _a[117] ), .Z( _aa[58] ) );
XOR2UD1BWP30P140 U59 ( .A1( _a[118] ), .A2( _a[119] ), .Z( _aa[59] ) );
XOR2UD1BWP30P140 U60 ( .A1( _a[120] ), .A2( _a[121] ), .Z( _aa[60] ) );
XOR2UD1BWP30P140 U61 ( .A1( _a[122] ), .A2( _a[123] ), .Z( _aa[61] ) );
XOR2UD1BWP30P140 U62 ( .A1( _a[124] ), .A2( _a[125] ), .Z( _aa[62] ) );
XOR2UD1BWP30P140 U63 ( .A1( _a[126] ), .A2( _a[127] ), .Z( _aa[63] ) );
XOR2UD1BWP30P140 U64 ( .A1( _b[0] ), .A2( _b[1] ), .Z( _bb[0] ) );
XOR2UD1BWP30P140 U65 ( .A1( _b[2] ), .A2( _b[3] ), .Z( _bb[1] ) );
XOR2UD1BWP30P140 U66 ( .A1( _b[4] ), .A2( _b[5] ), .Z( _bb[2] ) );
XOR2UD1BWP30P140 U67 ( .A1( _b[6] ), .A2( _b[7] ), .Z( _bb[3] ) );
XOR2UD1BWP30P140 U68 ( .A1( _b[8] ), .A2( _b[9] ), .Z( _bb[4] ) );
XOR2UD1BWP30P140 U69 ( .A1( _b[10] ), .A2( _b[11] ), .Z( _bb[5] ) );
XOR2UD1BWP30P140 U70 ( .A1( _b[12] ), .A2( _b[13] ), .Z( _bb[6] ) );
XOR2UD1BWP30P140 U71 ( .A1( _b[14] ), .A2( _b[15] ), .Z( _bb[7] ) );
XOR2UD1BWP30P140 U72 ( .A1( _b[16] ), .A2( _b[17] ), .Z( _bb[8] ) );
XOR2UD1BWP30P140 U73 ( .A1( _b[18] ), .A2( _b[19] ), .Z( _bb[9] ) );
XOR2UD1BWP30P140 U74 ( .A1( _b[20] ), .A2( _b[21] ), .Z( _bb[10] ) );
XOR2UD1BWP30P140 U75 ( .A1( _b[22] ), .A2( _b[23] ), .Z( _bb[11] ) );
XOR2UD1BWP30P140 U76 ( .A1( _b[24] ), .A2( _b[25] ), .Z( _bb[12] ) );
XOR2UD1BWP30P140 U77 ( .A1( _b[26] ), .A2( _b[27] ), .Z( _bb[13] ) );
XOR2UD1BWP30P140 U78 ( .A1( _b[28] ), .A2( _b[29] ), .Z( _bb[14] ) );
XOR2UD1BWP30P140 U79 ( .A1( _b[30] ), .A2( _b[31] ), .Z( _bb[15] ) );
XOR2UD1BWP30P140 U80 ( .A1( _b[32] ), .A2( _b[33] ), .Z( _bb[16] ) );
XOR2UD1BWP30P140 U81 ( .A1( _b[34] ), .A2( _b[35] ), .Z( _bb[17] ) );
XOR2UD1BWP30P140 U82 ( .A1( _b[36] ), .A2( _b[37] ), .Z( _bb[18] ) );
XOR2UD1BWP30P140 U83 ( .A1( _b[38] ), .A2( _b[39] ), .Z( _bb[19] ) );
XOR2UD1BWP30P140 U84 ( .A1( _b[40] ), .A2( _b[41] ), .Z( _bb[20] ) );
XOR2UD1BWP30P140 U85 ( .A1( _b[42] ), .A2( _b[43] ), .Z( _bb[21] ) );
XOR2UD1BWP30P140 U86 ( .A1( _b[44] ), .A2( _b[45] ), .Z( _bb[22] ) );
XOR2UD1BWP30P140 U87 ( .A1( _b[46] ), .A2( _b[47] ), .Z( _bb[23] ) );
XOR2UD1BWP30P140 U88 ( .A1( _b[48] ), .A2( _b[49] ), .Z( _bb[24] ) );
XOR2UD1BWP30P140 U89 ( .A1( _b[50] ), .A2( _b[51] ), .Z( _bb[25] ) );
XOR2UD1BWP30P140 U90 ( .A1( _b[52] ), .A2( _b[53] ), .Z( _bb[26] ) );
XOR2UD1BWP30P140 U91 ( .A1( _b[54] ), .A2( _b[55] ), .Z( _bb[27] ) );
XOR2UD1BWP30P140 U92 ( .A1( _b[56] ), .A2( _b[57] ), .Z( _bb[28] ) );
XOR2UD1BWP30P140 U93 ( .A1( _b[58] ), .A2( _b[59] ), .Z( _bb[29] ) );
XOR2UD1BWP30P140 U94 ( .A1( _b[60] ), .A2( _b[61] ), .Z( _bb[30] ) );
XOR2UD1BWP30P140 U95 ( .A1( _b[62] ), .A2( _b[63] ), .Z( _bb[31] ) );
XOR2UD1BWP30P140 U96 ( .A1( _b[64] ), .A2( _b[65] ), .Z( _bb[32] ) );
XOR2UD1BWP30P140 U97 ( .A1( _b[66] ), .A2( _b[67] ), .Z( _bb[33] ) );
XOR2UD1BWP30P140 U98 ( .A1( _b[68] ), .A2( _b[69] ), .Z( _bb[34] ) );
XOR2UD1BWP30P140 U99 ( .A1( _b[70] ), .A2( _b[71] ), .Z( _bb[35] ) );
XOR2UD1BWP30P140 U100 ( .A1( _b[72] ), .A2( _b[73] ), .Z( _bb[36] ) );
XOR2UD1BWP30P140 U101 ( .A1( _b[74] ), .A2( _b[75] ), .Z( _bb[37] ) );
XOR2UD1BWP30P140 U102 ( .A1( _b[76] ), .A2( _b[77] ), .Z( _bb[38] ) );
XOR2UD1BWP30P140 U103 ( .A1( _b[78] ), .A2( _b[79] ), .Z( _bb[39] ) );
XOR2UD1BWP30P140 U104 ( .A1( _b[80] ), .A2( _b[81] ), .Z( _bb[40] ) );
XOR2UD1BWP30P140 U105 ( .A1( _b[82] ), .A2( _b[83] ), .Z( _bb[41] ) );
XOR2UD1BWP30P140 U106 ( .A1( _b[84] ), .A2( _b[85] ), .Z( _bb[42] ) );
XOR2UD1BWP30P140 U107 ( .A1( _b[86] ), .A2( _b[87] ), .Z( _bb[43] ) );
XOR2UD1BWP30P140 U108 ( .A1( _b[88] ), .A2( _b[89] ), .Z( _bb[44] ) );
XOR2UD1BWP30P140 U109 ( .A1( _b[90] ), .A2( _b[91] ), .Z( _bb[45] ) );
XOR2UD1BWP30P140 U110 ( .A1( _b[92] ), .A2( _b[93] ), .Z( _bb[46] ) );
XOR2UD1BWP30P140 U111 ( .A1( _b[94] ), .A2( _b[95] ), .Z( _bb[47] ) );
XOR2UD1BWP30P140 U112 ( .A1( _b[96] ), .A2( _b[97] ), .Z( _bb[48] ) );
XOR2UD1BWP30P140 U113 ( .A1( _b[98] ), .A2( _b[99] ), .Z( _bb[49] ) );
XOR2UD1BWP30P140 U114 ( .A1( _b[100] ), .A2( _b[101] ), .Z( _bb[50] ) );
XOR2UD1BWP30P140 U115 ( .A1( _b[102] ), .A2( _b[103] ), .Z( _bb[51] ) );
XOR2UD1BWP30P140 U116 ( .A1( _b[104] ), .A2( _b[105] ), .Z( _bb[52] ) );
XOR2UD1BWP30P140 U117 ( .A1( _b[106] ), .A2( _b[107] ), .Z( _bb[53] ) );
XOR2UD1BWP30P140 U118 ( .A1( _b[108] ), .A2( _b[109] ), .Z( _bb[54] ) );
XOR2UD1BWP30P140 U119 ( .A1( _b[110] ), .A2( _b[111] ), .Z( _bb[55] ) );
XOR2UD1BWP30P140 U120 ( .A1( _b[112] ), .A2( _b[113] ), .Z( _bb[56] ) );
XOR2UD1BWP30P140 U121 ( .A1( _b[114] ), .A2( _b[115] ), .Z( _bb[57] ) );
XOR2UD1BWP30P140 U122 ( .A1( _b[116] ), .A2( _b[117] ), .Z( _bb[58] ) );
XOR2UD1BWP30P140 U123 ( .A1( _b[118] ), .A2( _b[119] ), .Z( _bb[59] ) );
XOR2UD1BWP30P140 U124 ( .A1( _b[120] ), .A2( _b[121] ), .Z( _bb[60] ) );
XOR2UD1BWP30P140 U125 ( .A1( _b[122] ), .A2( _b[123] ), .Z( _bb[61] ) );
XOR2UD1BWP30P140 U126 ( .A1( _b[124] ), .A2( _b[125] ), .Z( _bb[62] ) );
XOR2UD1BWP30P140 U127 ( .A1( _b[126] ), .A2( _b[127] ), .Z( _bb[63] ) );
endmodule
