module OKA_8bit_0_19 ( a, b, y );
input [7:0] a;
input [7:0] b;
output [7:0] y;
wire [7:0] _a;
wire [7:0] _b;
wire [7:0] _y;
wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;
assign _a = a;
assign _b = b;
assign y = _y;
XOR2UD1BWP30P140 U1 ( .A1( n84 ), .A2( n83 ), .Z( _y[7] ) );
XOR4D1BWP30P140 U2 ( .A1( n78 ), .A2( n77 ), .A3( n76 ), .A4( n75 ), .Z( n84 ) );
XOR4D1BWP30P140 U3 ( .A1( n82 ), .A2( n81 ), .A3( n80 ), .A4( n79 ), .Z( n83 ) );
CKND2D1BWP30P140 U4 ( .A1( _b[5] ), .A2( _a[2] ), .ZN( n78 ) );
XOR4D1BWP30P140 U5 ( .A1( n66 ), .A2( n65 ), .A3( n64 ), .A4( n63 ), .Z( _y[5] ) );
CKND2D1BWP30P140 U6 ( .A1( _b[0] ), .A2( _a[5] ), .ZN( n63 ) );
NR2D1BWP30P140 U7 ( .A1( n87 ), .A2( n86 ), .ZN( n66 ) );
NR2D1BWP30P140 U8 ( .A1( n88 ), .A2( n85 ), .ZN( n65 ) );
XOR4D1BWP30P140 U9 ( .A1( n70 ), .A2( n69 ), .A3( n68 ), .A4( n67 ), .Z( n74 ) );
CKND2D1BWP30P140 U10 ( .A1( _b[4] ), .A2( _a[2] ), .ZN( n70 ) );
CKND2D1BWP30P140 U11 ( .A1( _a[0] ), .A2( _b[6] ), .ZN( n67 ) );
CKND2D1BWP30P140 U12 ( .A1( _b[3] ), .A2( _a[3] ), .ZN( n69 ) );
XOR3UD1BWP30P140 U13 ( .A1( n59 ), .A2( n58 ), .A3( n57 ), .Z( _y[4] ) );
CKND2D1BWP30P140 U14 ( .A1( _b[0] ), .A2( _a[4] ), .ZN( n58 ) );
NR2D1BWP30P140 U15 ( .A1( n87 ), .A2( n85 ), .ZN( n59 ) );
XOR3UD1BWP30P140 U16 ( .A1( n56 ), .A2( n55 ), .A3( n54 ), .Z( n57 ) );
XOR3UD1BWP30P140 U17 ( .A1( n49 ), .A2( n48 ), .A3( n47 ), .Z( _y[2] ) );
AN2D1BWP30P140 U18 ( .A1( _a[2] ), .A2( _b[0] ), .Z( n47 ) );
AN2D1BWP30P140 U19 ( .A1( _a[0] ), .A2( _b[2] ), .Z( n48 ) );
INR2D1BWP30P140 U20 ( .A1( _a[1] ), .B1( n85 ), .ZN( n49 ) );
INVD1BWP30P140 U21 ( .I( _b[2] ), .ZN( n86 ) );
AN2D1BWP30P140 U22 ( .A1( _a[0] ), .A2( _b[0] ), .Z( _y[0] ) );
XOR3UD1BWP30P140 U23 ( .A1( n62 ), .A2( n61 ), .A3( n60 ), .Z( n64 ) );
CKND2D1BWP30P140 U24 ( .A1( _b[3] ), .A2( _a[2] ), .ZN( n60 ) );
CKND2D1BWP30P140 U25 ( .A1( _b[4] ), .A2( _a[1] ), .ZN( n61 ) );
CKND2D1BWP30P140 U26 ( .A1( _b[5] ), .A2( _a[0] ), .ZN( n62 ) );
CKND2D1BWP30P140 U27 ( .A1( _b[3] ), .A2( _a[1] ), .ZN( n55 ) );
CKND2D1BWP30P140 U28 ( .A1( _b[7] ), .A2( _a[0] ), .ZN( n75 ) );
INVD1BWP30P140 U29 ( .I( _a[4] ), .ZN( n88 ) );
INVD1BWP30P140 U30 ( .I( _a[3] ), .ZN( n87 ) );
CKND2D1BWP30P140 U31 ( .A1( _b[2] ), .A2( _a[5] ), .ZN( n79 ) );
CKND2D1BWP30P140 U32 ( .A1( _b[4] ), .A2( _a[0] ), .ZN( n56 ) );
CKND2D1BWP30P140 U33 ( .A1( _b[4] ), .A2( _a[3] ), .ZN( n77 ) );
CKND2D1BWP30P140 U34 ( .A1( _b[6] ), .A2( _a[1] ), .ZN( n76 ) );
CKND2D1BWP30P140 U35 ( .A1( _b[5] ), .A2( _a[1] ), .ZN( n68 ) );
CKND2D1BWP30P140 U36 ( .A1( _b[3] ), .A2( _a[4] ), .ZN( n80 ) );
CKND2D1BWP30P140 U37 ( .A1( _b[0] ), .A2( _a[7] ), .ZN( n81 ) );
CKND2D1BWP30P140 U38 ( .A1( _b[2] ), .A2( _a[2] ), .ZN( n54 ) );
CKND2D1BWP30P140 U39 ( .A1( _b[2] ), .A2( _a[1] ), .ZN( n51 ) );
XOR2UD1BWP30P140 U40 ( .A1( n46 ), .A2( n45 ), .Z( _y[1] ) );
CKND2D1BWP30P140 U41 ( .A1( _b[0] ), .A2( _a[1] ), .ZN( n46 ) );
CKND2D1BWP30P140 U42 ( .A1( _b[1] ), .A2( _a[0] ), .ZN( n45 ) );
INVD1BWP30P140 U43 ( .I( _b[1] ), .ZN( n85 ) );
XOR4D1BWP30P140 U44 ( .A1( n53 ), .A2( n52 ), .A3( n51 ), .A4( n50 ), .Z( _y[3] ) );
CKND2D1BWP30P140 U45 ( .A1( _b[3] ), .A2( _a[0] ), .ZN( n50 ) );
CKND2D1BWP30P140 U46 ( .A1( _b[1] ), .A2( _a[2] ), .ZN( n53 ) );
CKND2D1BWP30P140 U47 ( .A1( _b[0] ), .A2( _a[3] ), .ZN( n52 ) );
XOR4D1BWP30P140 U48 ( .A1( n74 ), .A2( n73 ), .A3( n72 ), .A4( n71 ), .Z( _y[6] ) );
CKND2D1BWP30P140 U49 ( .A1( _b[0] ), .A2( _a[6] ), .ZN( n71 ) );
CKND2D1BWP30P140 U50 ( .A1( _b[1] ), .A2( _a[5] ), .ZN( n72 ) );
NR2D1BWP30P140 U51 ( .A1( n88 ), .A2( n86 ), .ZN( n73 ) );
CKND2D1BWP30P140 U52 ( .A1( _b[1] ), .A2( _a[6] ), .ZN( n82 ) );
endmodule
