module OKA_16bit_15 ( a, b, y );
input [15:0] a;
input [15:0] b;
output [30:0] y;
wire [30:0] _y;
wire [7:0] aa;
wire [7:0] bb;
wire [7:0] al;
wire [7:0] ah;
wire [7:0] bl;
wire [7:0] bh;
wire [14:0] z1;
wire [6:0] o;
assign al = a[7:0];
assign ah = a[15:8];
assign bl = b[7:0];
assign bh = b[15:8];
assign y = _y;
s_16bit_15 s16_u ( .a( { ah, al } ), .b( { bh, bl } ), .aa( aa ), .bb( bb ) );
OKA_8bit_0_15 mul8_0 ( .a( al ), .b( bl ), .y( _y[7:0] ) );
OKA_8bit_1_15 mul8_1 ( .a( aa ), .b( bb ), .y( z1 ) );
OKA_8bit_2_15 mul8_2 ( .a( ah ), .b( bh ), .y( _y[30:23] ) );
OS_XOR2_15 os_xor2_u ( .a0( al ), .b0( bl ), .a1( ah ), .b1( bh ), .y( o ) );
os_16bit_15 os16_u ( .z0( _y[7:0] ), .z1( z1 ), .z2( _y[30:23] ), .o( o ), .y( _y[22:8] ) );
endmodule
