module OS_XOR2_17 ( a0, b0, a1, b1, y );
input [7:0] a0;
input [7:0] b0;
input [7:0] a1;
input [7:0] b1;
output [6:0] y;
wire [7:0] _a0;
wire [7:0] _b0;
wire [7:0] _a1;
wire [7:0] _b1;
wire [6:0] _y;
wire n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140;
assign _a0 = a0;
assign _b0 = b0;
assign _a1 = a1;
assign _b1 = b1;
assign y = _y;
XOR2UD1BWP30P140 U1 ( .A1( n90 ), .A2( n89 ), .Z( _y[1] ) );
XOR4D1BWP30P140 U2 ( .A1( n84 ), .A2( n83 ), .A3( n82 ), .A4( n81 ), .Z( n90 ) );
XOR4D1BWP30P140 U3 ( .A1( n88 ), .A2( n87 ), .A3( n86 ), .A4( n85 ), .Z( n89 ) );
CKND2D1BWP30P140 U4 ( .A1( _a0[4] ), .A2( _b0[5] ), .ZN( n84 ) );
XOR2UD1BWP30P140 U5 ( .A1( n80 ), .A2( n79 ), .Z( _y[0] ) );
XOR4D1BWP30P140 U6 ( .A1( n74 ), .A2( n73 ), .A3( n72 ), .A4( n71 ), .Z( n80 ) );
XOR4D1BWP30P140 U7 ( .A1( n78 ), .A2( n77 ), .A3( n76 ), .A4( n75 ), .Z( n79 ) );
CKND2D1BWP30P140 U8 ( .A1( _a0[3] ), .A2( _b0[5] ), .ZN( n74 ) );
XOR2UD1BWP30P140 U9 ( .A1( n120 ), .A2( n119 ), .Z( _y[4] ) );
XOR4D1BWP30P140 U10 ( .A1( n114 ), .A2( n113 ), .A3( n112 ), .A4( n111 ), .Z( n120 ) );
XOR4D1BWP30P140 U11 ( .A1( n118 ), .A2( n117 ), .A3( n116 ), .A4( n115 ), .Z( n119 ) );
CKND2D1BWP30P140 U12 ( .A1( _b0[5] ), .A2( _a0[7] ), .ZN( n114 ) );
XOR2UD1BWP30P140 U13 ( .A1( n110 ), .A2( n109 ), .Z( _y[3] ) );
XOR4D1BWP30P140 U14 ( .A1( n104 ), .A2( n103 ), .A3( n102 ), .A4( n101 ), .Z( n110 ) );
XOR4D1BWP30P140 U15 ( .A1( n108 ), .A2( n107 ), .A3( n106 ), .A4( n105 ), .Z( n109 ) );
CKND2D1BWP30P140 U16 ( .A1( _b0[5] ), .A2( _a0[6] ), .ZN( n104 ) );
XOR2UD1BWP30P140 U17 ( .A1( n100 ), .A2( n99 ), .Z( _y[2] ) );
XOR4D1BWP30P140 U18 ( .A1( n94 ), .A2( n93 ), .A3( n92 ), .A4( n91 ), .Z( n100 ) );
XOR4D1BWP30P140 U19 ( .A1( n98 ), .A2( n97 ), .A3( n96 ), .A4( n95 ), .Z( n99 ) );
CKND2D1BWP30P140 U20 ( .A1( _b0[5] ), .A2( _a0[5] ), .ZN( n94 ) );
XOR2UD1BWP30P140 U21 ( .A1( n140 ), .A2( n139 ), .Z( _y[6] ) );
XOR4D1BWP30P140 U22 ( .A1( n134 ), .A2( n133 ), .A3( n132 ), .A4( n131 ), .Z( n140 ) );
XOR4D1BWP30P140 U23 ( .A1( n138 ), .A2( n137 ), .A3( n136 ), .A4( n135 ), .Z( n139 ) );
CKND2D1BWP30P140 U24 ( .A1( _b1[5] ), .A2( _a1[1] ), .ZN( n134 ) );
XOR2UD1BWP30P140 U25 ( .A1( n130 ), .A2( n129 ), .Z( _y[5] ) );
XOR4D1BWP30P140 U26 ( .A1( n124 ), .A2( n123 ), .A3( n122 ), .A4( n121 ), .Z( n130 ) );
XOR4D1BWP30P140 U27 ( .A1( n128 ), .A2( n127 ), .A3( n126 ), .A4( n125 ), .Z( n129 ) );
CKND2D1BWP30P140 U28 ( .A1( _b1[5] ), .A2( _a1[0] ), .ZN( n124 ) );
CKND2D1BWP30P140 U29 ( .A1( _b1[1] ), .A2( _a1[1] ), .ZN( n98 ) );
CKND2D1BWP30P140 U30 ( .A1( _b1[1] ), .A2( _a1[0] ), .ZN( n88 ) );
CKND2D1BWP30P140 U31 ( .A1( _a0[6] ), .A2( _b0[7] ), .ZN( n121 ) );
CKND2D1BWP30P140 U32 ( .A1( _a0[5] ), .A2( _b0[7] ), .ZN( n111 ) );
CKND2D1BWP30P140 U33 ( .A1( _b1[2] ), .A2( _a1[1] ), .ZN( n105 ) );
CKND2D1BWP30P140 U34 ( .A1( _a0[4] ), .A2( _b0[7] ), .ZN( n101 ) );
CKND2D1BWP30P140 U35 ( .A1( _a0[3] ), .A2( _b0[7] ), .ZN( n91 ) );
CKND2D1BWP30P140 U36 ( .A1( _a0[2] ), .A2( _b0[7] ), .ZN( n81 ) );
CKND2D1BWP30P140 U37 ( .A1( _b0[2] ), .A2( _a0[6] ), .ZN( n75 ) );
CKND2D1BWP30P140 U38 ( .A1( _a0[1] ), .A2( _b0[7] ), .ZN( n71 ) );
CKND2D1BWP30P140 U39 ( .A1( _b1[2] ), .A2( _a1[0] ), .ZN( n95 ) );
CKND2D1BWP30P140 U40 ( .A1( _b1[1] ), .A2( _a1[3] ), .ZN( n118 ) );
CKND2D1BWP30P140 U41 ( .A1( _b0[7] ), .A2( _a0[7] ), .ZN( n131 ) );
CKND2D1BWP30P140 U42 ( .A1( _b0[2] ), .A2( _a0[7] ), .ZN( n85 ) );
CKND2D1BWP30P140 U43 ( .A1( _b1[1] ), .A2( _a1[4] ), .ZN( n128 ) );
CKND2D1BWP30P140 U44 ( .A1( _b1[1] ), .A2( _a1[2] ), .ZN( n108 ) );
CKND2D1BWP30P140 U45 ( .A1( _b1[2] ), .A2( _a1[3] ), .ZN( n125 ) );
CKND2D1BWP30P140 U46 ( .A1( _b1[2] ), .A2( _a1[4] ), .ZN( n135 ) );
CKND2D1BWP30P140 U47 ( .A1( _b1[2] ), .A2( _a1[2] ), .ZN( n115 ) );
CKND2D1BWP30P140 U48 ( .A1( _b1[4] ), .A2( _a1[1] ), .ZN( n123 ) );
CKND2D1BWP30P140 U49 ( .A1( _b0[4] ), .A2( _a0[6] ), .ZN( n93 ) );
CKND2D1BWP30P140 U50 ( .A1( _b1[0] ), .A2( _a1[1] ), .ZN( n87 ) );
CKND2D1BWP30P140 U51 ( .A1( _b0[4] ), .A2( _a0[5] ), .ZN( n83 ) );
CKND2D1BWP30P140 U52 ( .A1( _b1[4] ), .A2( _a1[0] ), .ZN( n113 ) );
CKND2D1BWP30P140 U53 ( .A1( _b1[0] ), .A2( _a1[0] ), .ZN( n77 ) );
CKND2D1BWP30P140 U54 ( .A1( _b1[3] ), .A2( _a1[1] ), .ZN( n116 ) );
CKND2D1BWP30P140 U55 ( .A1( _a0[6] ), .A2( _b0[6] ), .ZN( n112 ) );
CKND2D1BWP30P140 U56 ( .A1( _a0[5] ), .A2( _b0[6] ), .ZN( n102 ) );
CKND2D1BWP30P140 U57 ( .A1( _a0[4] ), .A2( _b0[6] ), .ZN( n92 ) );
CKND2D1BWP30P140 U58 ( .A1( _b0[3] ), .A2( _a0[6] ), .ZN( n86 ) );
CKND2D1BWP30P140 U59 ( .A1( _a0[3] ), .A2( _b0[6] ), .ZN( n82 ) );
CKND2D1BWP30P140 U60 ( .A1( _b0[3] ), .A2( _a0[5] ), .ZN( n76 ) );
CKND2D1BWP30P140 U61 ( .A1( _a0[2] ), .A2( _b0[6] ), .ZN( n72 ) );
CKND2D1BWP30P140 U62 ( .A1( _b0[4] ), .A2( _a0[7] ), .ZN( n103 ) );
CKND2D1BWP30P140 U63 ( .A1( _b1[6] ), .A2( _a1[0] ), .ZN( n132 ) );
CKND2D1BWP30P140 U64 ( .A1( _b1[3] ), .A2( _a1[0] ), .ZN( n106 ) );
CKND2D1BWP30P140 U65 ( .A1( _b0[6] ), .A2( _a0[7] ), .ZN( n122 ) );
CKND2D1BWP30P140 U66 ( .A1( _b0[3] ), .A2( _a0[7] ), .ZN( n96 ) );
CKND2D1BWP30P140 U67 ( .A1( _b1[1] ), .A2( _a1[5] ), .ZN( n138 ) );
CKND2D1BWP30P140 U68 ( .A1( _b1[0] ), .A2( _a1[3] ), .ZN( n107 ) );
CKND2D1BWP30P140 U69 ( .A1( _b1[4] ), .A2( _a1[2] ), .ZN( n133 ) );
CKND2D1BWP30P140 U70 ( .A1( _b1[0] ), .A2( _a1[4] ), .ZN( n117 ) );
CKND2D1BWP30P140 U71 ( .A1( _b1[0] ), .A2( _a1[2] ), .ZN( n97 ) );
CKND2D1BWP30P140 U72 ( .A1( _b1[3] ), .A2( _a1[3] ), .ZN( n136 ) );
CKND2D1BWP30P140 U73 ( .A1( _b1[3] ), .A2( _a1[2] ), .ZN( n126 ) );
CKND2D1BWP30P140 U74 ( .A1( _b1[0] ), .A2( _a1[5] ), .ZN( n127 ) );
CKND2D1BWP30P140 U75 ( .A1( _b0[4] ), .A2( _a0[4] ), .ZN( n73 ) );
CKND2D1BWP30P140 U76 ( .A1( _b0[1] ), .A2( _a0[7] ), .ZN( n78 ) );
CKND2D1BWP30P140 U77 ( .A1( _b1[0] ), .A2( _a1[6] ), .ZN( n137 ) );
endmodule
