module OKA_8bit_2_20 ( a, b, y );
input [7:0] a;
input [7:0] b;
output [7:0] y;
wire [7:0] _a;
wire [7:0] _b;
wire [7:0] _y;
wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;
assign _a = a;
assign _b = b;
assign y = _y;
XOR2UD1BWP30P140 U1 ( .A1( n54 ), .A2( n53 ), .Z( _y[0] ) );
XOR4D1BWP30P140 U2 ( .A1( n48 ), .A2( n47 ), .A3( n46 ), .A4( n45 ), .Z( n54 ) );
XOR4D1BWP30P140 U3 ( .A1( n52 ), .A2( n51 ), .A3( n50 ), .A4( n49 ), .Z( n53 ) );
CKND2D1BWP30P140 U4 ( .A1( _a[2] ), .A2( _b[5] ), .ZN( n48 ) );
XOR4D1BWP30P140 U5 ( .A1( n79 ), .A2( n78 ), .A3( n77 ), .A4( n76 ), .Z( _y[4] ) );
CKND2D1BWP30P140 U6 ( .A1( _b[5] ), .A2( _a[6] ), .ZN( n79 ) );
CKND2D1BWP30P140 U7 ( .A1( _a[4] ), .A2( _b[7] ), .ZN( n76 ) );
CKND2D1BWP30P140 U8 ( .A1( _b[4] ), .A2( _a[7] ), .ZN( n78 ) );
XOR4D1BWP30P140 U9 ( .A1( n69 ), .A2( n68 ), .A3( n67 ), .A4( n66 ), .Z( _y[2] ) );
CKND2D1BWP30P140 U10 ( .A1( _b[2] ), .A2( _a[7] ), .ZN( n66 ) );
NR2D1BWP30P140 U11 ( .A1( n87 ), .A2( n86 ), .ZN( n69 ) );
NR2D1BWP30P140 U12 ( .A1( n88 ), .A2( n85 ), .ZN( n68 ) );
XOR4D1BWP30P140 U13 ( .A1( n62 ), .A2( n61 ), .A3( n60 ), .A4( n59 ), .Z( _y[1] ) );
CKND2D1BWP30P140 U14 ( .A1( _b[1] ), .A2( _a[7] ), .ZN( n59 ) );
CKND2D1BWP30P140 U15 ( .A1( _b[2] ), .A2( _a[6] ), .ZN( n60 ) );
NR2D1BWP30P140 U16 ( .A1( n87 ), .A2( n85 ), .ZN( n61 ) );
XOR4D1BWP30P140 U17 ( .A1( n58 ), .A2( n57 ), .A3( n56 ), .A4( n55 ), .Z( n62 ) );
CKND2D1BWP30P140 U18 ( .A1( _a[3] ), .A2( _b[5] ), .ZN( n58 ) );
CKND2D1BWP30P140 U19 ( .A1( _a[1] ), .A2( _b[7] ), .ZN( n55 ) );
CKND2D1BWP30P140 U20 ( .A1( _b[4] ), .A2( _a[4] ), .ZN( n57 ) );
INVD1BWP30P140 U21 ( .I( _a[6] ), .ZN( n88 ) );
AN2D1BWP30P140 U22 ( .A1( _a[7] ), .A2( _b[7] ), .Z( _y[7] ) );
INVD1BWP30P140 U23 ( .I( _b[4] ), .ZN( n86 ) );
INVD1BWP30P140 U24 ( .I( _b[3] ), .ZN( n85 ) );
XOR3UD1BWP30P140 U25 ( .A1( n75 ), .A2( n74 ), .A3( n73 ), .Z( _y[3] ) );
CKND2D1BWP30P140 U26 ( .A1( _b[3] ), .A2( _a[7] ), .ZN( n74 ) );
NR2D1BWP30P140 U27 ( .A1( n88 ), .A2( n86 ), .ZN( n75 ) );
XOR3UD1BWP30P140 U28 ( .A1( n72 ), .A2( n71 ), .A3( n70 ), .Z( n73 ) );
XOR3UD1BWP30P140 U29 ( .A1( n65 ), .A2( n64 ), .A3( n63 ), .Z( n67 ) );
CKND2D1BWP30P140 U30 ( .A1( _a[4] ), .A2( _b[5] ), .ZN( n63 ) );
CKND2D1BWP30P140 U31 ( .A1( _a[3] ), .A2( _b[6] ), .ZN( n64 ) );
CKND2D1BWP30P140 U32 ( .A1( _a[2] ), .A2( _b[7] ), .ZN( n65 ) );
CKND2D1BWP30P140 U33 ( .A1( _a[4] ), .A2( _b[6] ), .ZN( n71 ) );
CKND2D1BWP30P140 U34 ( .A1( _b[1] ), .A2( _a[6] ), .ZN( n52 ) );
XOR2UD1BWP30P140 U35 ( .A1( n84 ), .A2( n83 ), .Z( _y[6] ) );
CKND2D1BWP30P140 U36 ( .A1( _b[6] ), .A2( _a[7] ), .ZN( n84 ) );
CKND2D1BWP30P140 U37 ( .A1( _a[6] ), .A2( _b[7] ), .ZN( n83 ) );
CKND2D1BWP30P140 U38 ( .A1( _a[0] ), .A2( _b[7] ), .ZN( n45 ) );
CKND2D1BWP30P140 U39 ( .A1( _b[2] ), .A2( _a[5] ), .ZN( n49 ) );
INVD1BWP30P140 U40 ( .I( _a[5] ), .ZN( n87 ) );
XOR3UD1BWP30P140 U41 ( .A1( n82 ), .A2( n81 ), .A3( n80 ), .Z( _y[5] ) );
AN2D1BWP30P140 U42 ( .A1( _a[7] ), .A2( _b[5] ), .Z( n80 ) );
AN2D1BWP30P140 U43 ( .A1( _b[7] ), .A2( _a[5] ), .Z( n81 ) );
INR2D1BWP30P140 U44 ( .A1( _b[6] ), .B1( n88 ), .ZN( n82 ) );
CKND2D1BWP30P140 U45 ( .A1( _a[3] ), .A2( _b[7] ), .ZN( n72 ) );
CKND2D1BWP30P140 U46 ( .A1( _a[3] ), .A2( _b[4] ), .ZN( n47 ) );
CKND2D1BWP30P140 U47 ( .A1( _b[0] ), .A2( _a[7] ), .ZN( n51 ) );
CKND2D1BWP30P140 U48 ( .A1( _a[1] ), .A2( _b[6] ), .ZN( n46 ) );
CKND2D1BWP30P140 U49 ( .A1( _a[2] ), .A2( _b[6] ), .ZN( n56 ) );
CKND2D1BWP30P140 U50 ( .A1( _a[5] ), .A2( _b[5] ), .ZN( n70 ) );
CKND2D1BWP30P140 U51 ( .A1( _b[3] ), .A2( _a[4] ), .ZN( n50 ) );
CKND2D1BWP30P140 U52 ( .A1( _a[5] ), .A2( _b[6] ), .ZN( n77 ) );
endmodule
