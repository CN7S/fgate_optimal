module OKA_8bit_1_20 ( a, b, y );
input [7:0] a;
input [7:0] b;
output [14:0] y;
wire [7:0] _a;
wire [7:0] _b;
wire [14:0] _y;
wire n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156;
assign _a = a;
assign _b = b;
assign y = _y;
INVD1BWP30P140 U1 ( .I( _a[6] ), .ZN( n156 ) );
INVD1BWP30P140 U2 ( .I( _b[3] ), .ZN( n151 ) );
INVD1BWP30P140 U3 ( .I( _b[2] ), .ZN( n150 ) );
INVD1BWP30P140 U4 ( .I( _b[4] ), .ZN( n152 ) );
XOR2UD1BWP30P140 U5 ( .A1( n93 ), .A2( n92 ), .Z( _y[13] ) );
CKND2D1BWP30P140 U6 ( .A1( _a[6] ), .A2( _b[7] ), .ZN( n92 ) );
CKND2D1BWP30P140 U7 ( .A1( _a[7] ), .A2( _b[6] ), .ZN( n93 ) );
INVD1BWP30P140 U8 ( .I( _a[3] ), .ZN( n153 ) );
CKND2D1BWP30P140 U9 ( .A1( _a[2] ), .A2( _b[5] ), .ZN( n127 ) );
INVD1BWP30P140 U10 ( .I( _a[4] ), .ZN( n154 ) );
CKND2D1BWP30P140 U11 ( .A1( _b[6] ), .A2( _a[4] ), .ZN( n80 ) );
CKND2D1BWP30P140 U12 ( .A1( _a[2] ), .A2( _b[6] ), .ZN( n135 ) );
CKND2D1BWP30P140 U13 ( .A1( _a[1] ), .A2( _b[6] ), .ZN( n125 ) );
CKND2D1BWP30P140 U14 ( .A1( _a[5] ), .A2( _b[6] ), .ZN( n86 ) );
CKND2D1BWP30P140 U15 ( .A1( _a[1] ), .A2( _b[3] ), .ZN( n104 ) );
CKND2D1BWP30P140 U16 ( .A1( _b[2] ), .A2( _a[2] ), .ZN( n103 ) );
INVD1BWP30P140 U17 ( .I( _a[5] ), .ZN( n155 ) );
CKND2D1BWP30P140 U18 ( .A1( _a[5] ), .A2( _b[5] ), .ZN( n79 ) );
CKND2D1BWP30P140 U19 ( .A1( _a[0] ), .A2( _b[7] ), .ZN( n124 ) );
CKND2D1BWP30P140 U20 ( .A1( _a[1] ), .A2( _b[5] ), .ZN( n117 ) );
CKND2D1BWP30P140 U21 ( .A1( _a[0] ), .A2( _b[4] ), .ZN( n105 ) );
CKND2D1BWP30P140 U22 ( .A1( _b[7] ), .A2( _a[3] ), .ZN( n81 ) );
CKND2D1BWP30P140 U23 ( .A1( _b[4] ), .A2( _a[3] ), .ZN( n126 ) );
CKND2D1BWP30P140 U24 ( .A1( _b[0] ), .A2( _a[7] ), .ZN( n130 ) );
CKND2D1BWP30P140 U25 ( .A1( _b[3] ), .A2( _a[4] ), .ZN( n129 ) );
CKND2D1BWP30P140 U26 ( .A1( _a[1] ), .A2( _b[2] ), .ZN( n100 ) );
CKND2D1BWP30P140 U27 ( .A1( _a[5] ), .A2( _b[2] ), .ZN( n128 ) );
XOR4D1BWP30P140 U28 ( .A1( n137 ), .A2( n136 ), .A3( n135 ), .A4( n134 ), .Z( n141 ) );
CKND2D1BWP30P140 U29 ( .A1( _a[3] ), .A2( _b[5] ), .ZN( n137 ) );
CKND2D1BWP30P140 U30 ( .A1( _a[1] ), .A2( _b[7] ), .ZN( n134 ) );
CKND2D1BWP30P140 U31 ( .A1( _b[4] ), .A2( _a[4] ), .ZN( n136 ) );
XOR4D1BWP30P140 U32 ( .A1( n119 ), .A2( n118 ), .A3( n117 ), .A4( n116 ), .Z( n123 ) );
CKND2D1BWP30P140 U33 ( .A1( _b[4] ), .A2( _a[2] ), .ZN( n119 ) );
CKND2D1BWP30P140 U34 ( .A1( _b[3] ), .A2( _a[3] ), .ZN( n118 ) );
CKND2D1BWP30P140 U35 ( .A1( _a[0] ), .A2( _b[6] ), .ZN( n116 ) );
XOR4D1BWP30P140 U36 ( .A1( n115 ), .A2( n114 ), .A3( n113 ), .A4( n112 ), .Z( _y[5] ) );
CKND2D1BWP30P140 U37 ( .A1( _b[0] ), .A2( _a[5] ), .ZN( n112 ) );
NR2D1BWP30P140 U38 ( .A1( n153 ), .A2( n150 ), .ZN( n115 ) );
NR2D1BWP30P140 U39 ( .A1( n154 ), .A2( n149 ), .ZN( n114 ) );
XOR4D1BWP30P140 U40 ( .A1( n148 ), .A2( n147 ), .A3( n146 ), .A4( n145 ), .Z( _y[9] ) );
CKND2D1BWP30P140 U41 ( .A1( _b[2] ), .A2( _a[7] ), .ZN( n145 ) );
NR2D1BWP30P140 U42 ( .A1( n155 ), .A2( n152 ), .ZN( n148 ) );
NR2D1BWP30P140 U43 ( .A1( n156 ), .A2( n151 ), .ZN( n147 ) );
XOR4D1BWP30P140 U44 ( .A1( n88 ), .A2( n87 ), .A3( n86 ), .A4( n85 ), .Z( _y[11] ) );
CKND2D1BWP30P140 U45 ( .A1( _a[6] ), .A2( _b[5] ), .ZN( n88 ) );
CKND2D1BWP30P140 U46 ( .A1( _b[7] ), .A2( _a[4] ), .ZN( n85 ) );
CKND2D1BWP30P140 U47 ( .A1( _b[4] ), .A2( _a[7] ), .ZN( n87 ) );
AN2D1BWP30P140 U48 ( .A1( _a[0] ), .A2( _b[0] ), .Z( _y[0] ) );
AN2D1BWP30P140 U49 ( .A1( _b[7] ), .A2( _a[7] ), .Z( _y[14] ) );
XOR3UD1BWP30P140 U50 ( .A1( n108 ), .A2( n107 ), .A3( n106 ), .Z( _y[4] ) );
CKND2D1BWP30P140 U51 ( .A1( _b[0] ), .A2( _a[4] ), .ZN( n107 ) );
NR2D1BWP30P140 U52 ( .A1( n153 ), .A2( n149 ), .ZN( n108 ) );
XOR3UD1BWP30P140 U53 ( .A1( n105 ), .A2( n104 ), .A3( n103 ), .Z( n106 ) );
XOR3UD1BWP30P140 U54 ( .A1( n84 ), .A2( n83 ), .A3( n82 ), .Z( _y[10] ) );
CKND2D1BWP30P140 U55 ( .A1( _b[3] ), .A2( _a[7] ), .ZN( n83 ) );
NR2D1BWP30P140 U56 ( .A1( n152 ), .A2( n156 ), .ZN( n84 ) );
XOR3UD1BWP30P140 U57 ( .A1( n81 ), .A2( n80 ), .A3( n79 ), .Z( n82 ) );
XOR3UD1BWP30P140 U58 ( .A1( n111 ), .A2( n110 ), .A3( n109 ), .Z( n113 ) );
CKND2D1BWP30P140 U59 ( .A1( _b[3] ), .A2( _a[2] ), .ZN( n109 ) );
CKND2D1BWP30P140 U60 ( .A1( _a[1] ), .A2( _b[4] ), .ZN( n110 ) );
CKND2D1BWP30P140 U61 ( .A1( _a[0] ), .A2( _b[5] ), .ZN( n111 ) );
XOR3UD1BWP30P140 U62 ( .A1( n144 ), .A2( n143 ), .A3( n142 ), .Z( n146 ) );
CKND2D1BWP30P140 U63 ( .A1( _b[5] ), .A2( _a[4] ), .ZN( n142 ) );
CKND2D1BWP30P140 U64 ( .A1( _b[6] ), .A2( _a[3] ), .ZN( n143 ) );
CKND2D1BWP30P140 U65 ( .A1( _b[7] ), .A2( _a[2] ), .ZN( n144 ) );
XOR3UD1BWP30P140 U66 ( .A1( n91 ), .A2( n90 ), .A3( n89 ), .Z( _y[12] ) );
AN2D1BWP30P140 U67 ( .A1( _b[5] ), .A2( _a[7] ), .Z( n89 ) );
AN2D1BWP30P140 U68 ( .A1( _b[7] ), .A2( _a[5] ), .Z( n90 ) );
INR2D1BWP30P140 U69 ( .A1( _b[6] ), .B1( n156 ), .ZN( n91 ) );
XOR3UD1BWP30P140 U70 ( .A1( n98 ), .A2( n97 ), .A3( n96 ), .Z( _y[2] ) );
AN2D1BWP30P140 U71 ( .A1( _a[2] ), .A2( _b[0] ), .Z( n96 ) );
AN2D1BWP30P140 U72 ( .A1( _a[0] ), .A2( _b[2] ), .Z( n97 ) );
INR2D1BWP30P140 U73 ( .A1( _a[1] ), .B1( n149 ), .ZN( n98 ) );
INVD1BWP30P140 U74 ( .I( _b[1] ), .ZN( n149 ) );
XOR2UD1BWP30P140 U75 ( .A1( n133 ), .A2( n132 ), .Z( _y[7] ) );
XOR4D1BWP30P140 U76 ( .A1( n131 ), .A2( n130 ), .A3( n129 ), .A4( n128 ), .Z( n132 ) );
XOR4D1BWP30P140 U77 ( .A1( n127 ), .A2( n126 ), .A3( n125 ), .A4( n124 ), .Z( n133 ) );
CKND2D1BWP30P140 U78 ( .A1( _b[1] ), .A2( _a[6] ), .ZN( n131 ) );
XOR2UD1BWP30P140 U79 ( .A1( n95 ), .A2( n94 ), .Z( _y[1] ) );
CKND2D1BWP30P140 U80 ( .A1( _b[0] ), .A2( _a[1] ), .ZN( n95 ) );
CKND2D1BWP30P140 U81 ( .A1( _a[0] ), .A2( _b[1] ), .ZN( n94 ) );
XOR4D1BWP30P140 U82 ( .A1( n141 ), .A2( n140 ), .A3( n139 ), .A4( n138 ), .Z( _y[8] ) );
CKND2D1BWP30P140 U83 ( .A1( _b[1] ), .A2( _a[7] ), .ZN( n138 ) );
CKND2D1BWP30P140 U84 ( .A1( _a[6] ), .A2( _b[2] ), .ZN( n139 ) );
NR2D1BWP30P140 U85 ( .A1( n155 ), .A2( n151 ), .ZN( n140 ) );
XOR4D1BWP30P140 U86 ( .A1( n123 ), .A2( n122 ), .A3( n121 ), .A4( n120 ), .Z( _y[6] ) );
CKND2D1BWP30P140 U87 ( .A1( _b[0] ), .A2( _a[6] ), .ZN( n120 ) );
CKND2D1BWP30P140 U88 ( .A1( _b[1] ), .A2( _a[5] ), .ZN( n121 ) );
NR2D1BWP30P140 U89 ( .A1( n154 ), .A2( n150 ), .ZN( n122 ) );
XOR4D1BWP30P140 U90 ( .A1( n102 ), .A2( n101 ), .A3( n100 ), .A4( n99 ), .Z( _y[3] ) );
CKND2D1BWP30P140 U91 ( .A1( _b[1] ), .A2( _a[2] ), .ZN( n102 ) );
CKND2D1BWP30P140 U92 ( .A1( _a[0] ), .A2( _b[3] ), .ZN( n99 ) );
CKND2D1BWP30P140 U93 ( .A1( _b[0] ), .A2( _a[3] ), .ZN( n101 ) );
endmodule
