module s_32bit_1 ( a, b, aa, bb );
input [31:0] a;
input [31:0] b;
output [15:0] aa;
output [15:0] bb;
wire [31:0] _a;
wire [31:0] _b;
wire [15:0] _aa;
wire [15:0] _bb;
assign _a = a;
assign _b = b;
assign aa = _aa;
assign bb = _bb;
XOR2UD1BWP30P140 U0 ( .A1( _a[0] ), .A2( _a[16] ), .Z( _aa[0] ) );
XOR2UD1BWP30P140 U1 ( .A1( _a[1] ), .A2( _a[17] ), .Z( _aa[1] ) );
XOR2UD1BWP30P140 U2 ( .A1( _a[2] ), .A2( _a[18] ), .Z( _aa[2] ) );
XOR2UD1BWP30P140 U3 ( .A1( _a[3] ), .A2( _a[19] ), .Z( _aa[3] ) );
XOR2UD1BWP30P140 U4 ( .A1( _a[4] ), .A2( _a[20] ), .Z( _aa[4] ) );
XOR2UD1BWP30P140 U5 ( .A1( _a[5] ), .A2( _a[21] ), .Z( _aa[5] ) );
XOR2UD1BWP30P140 U6 ( .A1( _a[6] ), .A2( _a[22] ), .Z( _aa[6] ) );
XOR2UD1BWP30P140 U7 ( .A1( _a[7] ), .A2( _a[23] ), .Z( _aa[7] ) );
XOR2UD1BWP30P140 U8 ( .A1( _a[8] ), .A2( _a[24] ), .Z( _aa[8] ) );
XOR2UD1BWP30P140 U9 ( .A1( _a[9] ), .A2( _a[25] ), .Z( _aa[9] ) );
XOR2UD1BWP30P140 U10 ( .A1( _a[10] ), .A2( _a[26] ), .Z( _aa[10] ) );
XOR2UD1BWP30P140 U11 ( .A1( _a[11] ), .A2( _a[27] ), .Z( _aa[11] ) );
XOR2UD1BWP30P140 U12 ( .A1( _a[12] ), .A2( _a[28] ), .Z( _aa[12] ) );
XOR2UD1BWP30P140 U13 ( .A1( _a[13] ), .A2( _a[29] ), .Z( _aa[13] ) );
XOR2UD1BWP30P140 U14 ( .A1( _a[14] ), .A2( _a[30] ), .Z( _aa[14] ) );
XOR2UD1BWP30P140 U15 ( .A1( _a[15] ), .A2( _a[31] ), .Z( _aa[15] ) );
XOR2UD1BWP30P140 U16 ( .A1( _b[0] ), .A2( _b[16] ), .Z( _bb[0] ) );
XOR2UD1BWP30P140 U17 ( .A1( _b[1] ), .A2( _b[17] ), .Z( _bb[1] ) );
XOR2UD1BWP30P140 U18 ( .A1( _b[2] ), .A2( _b[18] ), .Z( _bb[2] ) );
XOR2UD1BWP30P140 U19 ( .A1( _b[3] ), .A2( _b[19] ), .Z( _bb[3] ) );
XOR2UD1BWP30P140 U20 ( .A1( _b[4] ), .A2( _b[20] ), .Z( _bb[4] ) );
XOR2UD1BWP30P140 U21 ( .A1( _b[5] ), .A2( _b[21] ), .Z( _bb[5] ) );
XOR2UD1BWP30P140 U22 ( .A1( _b[6] ), .A2( _b[22] ), .Z( _bb[6] ) );
XOR2UD1BWP30P140 U23 ( .A1( _b[7] ), .A2( _b[23] ), .Z( _bb[7] ) );
XOR2UD1BWP30P140 U24 ( .A1( _b[8] ), .A2( _b[24] ), .Z( _bb[8] ) );
XOR2UD1BWP30P140 U25 ( .A1( _b[9] ), .A2( _b[25] ), .Z( _bb[9] ) );
XOR2UD1BWP30P140 U26 ( .A1( _b[10] ), .A2( _b[26] ), .Z( _bb[10] ) );
XOR2UD1BWP30P140 U27 ( .A1( _b[11] ), .A2( _b[27] ), .Z( _bb[11] ) );
XOR2UD1BWP30P140 U28 ( .A1( _b[12] ), .A2( _b[28] ), .Z( _bb[12] ) );
XOR2UD1BWP30P140 U29 ( .A1( _b[13] ), .A2( _b[29] ), .Z( _bb[13] ) );
XOR2UD1BWP30P140 U30 ( .A1( _b[14] ), .A2( _b[30] ), .Z( _bb[14] ) );
XOR2UD1BWP30P140 U31 ( .A1( _b[15] ), .A2( _b[31] ), .Z( _bb[15] ) );
endmodule
