module os_32bit_3 ( z0, z1, z2, y );
input [30:0] z0;
input [30:0] z1;
input [30:0] z2;
output [30:0] y;
wire [30:0] _z0;
wire [30:0] _z1;
wire [30:0] _z2;
wire [30:0] _y;
wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
assign _z0 = z0;
assign _z1 = z1;
assign _z2 = z2;
assign y = _y;
XOR2UD1BWP30P140 U0 ( .A1( _z2[0] ), .A2( _z0[16] ), .Z( n0 ) );
XOR2UD1BWP30P140 U1 ( .A1( _z2[1] ), .A2( _z0[17] ), .Z( n1 ) );
XOR2UD1BWP30P140 U2 ( .A1( _z2[2] ), .A2( _z0[18] ), .Z( n2 ) );
XOR2UD1BWP30P140 U3 ( .A1( _z2[3] ), .A2( _z0[19] ), .Z( n3 ) );
XOR2UD1BWP30P140 U4 ( .A1( _z2[4] ), .A2( _z0[20] ), .Z( n4 ) );
XOR2UD1BWP30P140 U5 ( .A1( _z2[5] ), .A2( _z0[21] ), .Z( n5 ) );
XOR2UD1BWP30P140 U6 ( .A1( _z2[6] ), .A2( _z0[22] ), .Z( n6 ) );
XOR2UD1BWP30P140 U7 ( .A1( _z2[7] ), .A2( _z0[23] ), .Z( n7 ) );
XOR2UD1BWP30P140 U8 ( .A1( _z2[8] ), .A2( _z0[24] ), .Z( n8 ) );
XOR2UD1BWP30P140 U9 ( .A1( _z2[9] ), .A2( _z0[25] ), .Z( n9 ) );
XOR2UD1BWP30P140 U10 ( .A1( _z2[10] ), .A2( _z0[26] ), .Z( n10 ) );
XOR2UD1BWP30P140 U11 ( .A1( _z2[11] ), .A2( _z0[27] ), .Z( n11 ) );
XOR2UD1BWP30P140 U12 ( .A1( _z2[12] ), .A2( _z0[28] ), .Z( n12 ) );
XOR2UD1BWP30P140 U13 ( .A1( _z2[13] ), .A2( _z0[29] ), .Z( n13 ) );
XOR2UD1BWP30P140 U14 ( .A1( _z2[14] ), .A2( _z0[30] ), .Z( n14 ) );
XOR3UD1BWP30P140 U15 ( .A1( _z1[0] ), .A2( _z0[0] ), .A3( n0 ), .Z( _y[0] ) );
XOR3UD1BWP30P140 U16 ( .A1( _z1[1] ), .A2( _z0[1] ), .A3( n1 ), .Z( _y[1] ) );
XOR3UD1BWP30P140 U17 ( .A1( _z1[2] ), .A2( _z0[2] ), .A3( n2 ), .Z( _y[2] ) );
XOR3UD1BWP30P140 U18 ( .A1( _z1[3] ), .A2( _z0[3] ), .A3( n3 ), .Z( _y[3] ) );
XOR3UD1BWP30P140 U19 ( .A1( _z1[4] ), .A2( _z0[4] ), .A3( n4 ), .Z( _y[4] ) );
XOR3UD1BWP30P140 U20 ( .A1( _z1[5] ), .A2( _z0[5] ), .A3( n5 ), .Z( _y[5] ) );
XOR3UD1BWP30P140 U21 ( .A1( _z1[6] ), .A2( _z0[6] ), .A3( n6 ), .Z( _y[6] ) );
XOR3UD1BWP30P140 U22 ( .A1( _z1[7] ), .A2( _z0[7] ), .A3( n7 ), .Z( _y[7] ) );
XOR3UD1BWP30P140 U23 ( .A1( _z1[8] ), .A2( _z0[8] ), .A3( n8 ), .Z( _y[8] ) );
XOR3UD1BWP30P140 U24 ( .A1( _z1[9] ), .A2( _z0[9] ), .A3( n9 ), .Z( _y[9] ) );
XOR3UD1BWP30P140 U25 ( .A1( _z1[10] ), .A2( _z0[10] ), .A3( n10 ), .Z( _y[10] ) );
XOR3UD1BWP30P140 U26 ( .A1( _z1[11] ), .A2( _z0[11] ), .A3( n11 ), .Z( _y[11] ) );
XOR3UD1BWP30P140 U27 ( .A1( _z1[12] ), .A2( _z0[12] ), .A3( n12 ), .Z( _y[12] ) );
XOR3UD1BWP30P140 U28 ( .A1( _z1[13] ), .A2( _z0[13] ), .A3( n13 ), .Z( _y[13] ) );
XOR3UD1BWP30P140 U29 ( .A1( _z1[14] ), .A2( _z0[14] ), .A3( n14 ), .Z( _y[14] ) );
XOR3UD1BWP30P140 U30 ( .A1( _z2[15] ), .A2( _z1[15] ), .A3( _z0[15] ), .Z( _y[15] ) );
XOR3UD1BWP30P140 U31 ( .A1( _z1[16] ), .A2( _z2[16] ), .A3( n0 ), .Z( _y[16] ) );
XOR3UD1BWP30P140 U32 ( .A1( _z1[17] ), .A2( _z2[17] ), .A3( n1 ), .Z( _y[17] ) );
XOR3UD1BWP30P140 U33 ( .A1( _z1[18] ), .A2( _z2[18] ), .A3( n2 ), .Z( _y[18] ) );
XOR3UD1BWP30P140 U34 ( .A1( _z1[19] ), .A2( _z2[19] ), .A3( n3 ), .Z( _y[19] ) );
XOR3UD1BWP30P140 U35 ( .A1( _z1[20] ), .A2( _z2[20] ), .A3( n4 ), .Z( _y[20] ) );
XOR3UD1BWP30P140 U36 ( .A1( _z1[21] ), .A2( _z2[21] ), .A3( n5 ), .Z( _y[21] ) );
XOR3UD1BWP30P140 U37 ( .A1( _z1[22] ), .A2( _z2[22] ), .A3( n6 ), .Z( _y[22] ) );
XOR3UD1BWP30P140 U38 ( .A1( _z1[23] ), .A2( _z2[23] ), .A3( n7 ), .Z( _y[23] ) );
XOR3UD1BWP30P140 U39 ( .A1( _z1[24] ), .A2( _z2[24] ), .A3( n8 ), .Z( _y[24] ) );
XOR3UD1BWP30P140 U40 ( .A1( _z1[25] ), .A2( _z2[25] ), .A3( n9 ), .Z( _y[25] ) );
XOR3UD1BWP30P140 U41 ( .A1( _z1[26] ), .A2( _z2[26] ), .A3( n10 ), .Z( _y[26] ) );
XOR3UD1BWP30P140 U42 ( .A1( _z1[27] ), .A2( _z2[27] ), .A3( n11 ), .Z( _y[27] ) );
XOR3UD1BWP30P140 U43 ( .A1( _z1[28] ), .A2( _z2[28] ), .A3( n12 ), .Z( _y[28] ) );
XOR3UD1BWP30P140 U44 ( .A1( _z1[29] ), .A2( _z2[29] ), .A3( n13 ), .Z( _y[29] ) );
XOR3UD1BWP30P140 U45 ( .A1( _z1[30] ), .A2( _z2[30] ), .A3( n14 ), .Z( _y[30] ) );
endmodule
