module s_16bit ( a, b, aa, bb );
input [15:0] a;
input [15:0] b;
output [7:0] aa;
output [7:0] bb;
wire [7:0] _aa;
wire [7:0] _bb;
wire [15:0] _a;
wire [15:0] _b;
assign _a = a;
assign _b = b;
assign aa = _aa;
assign bb = _bb;
XOR2UD1BWP30P140 U0 ( .A1( _a[0] ), .A2( _a[8] ), .Z( _aa[0] ) );
XOR2UD1BWP30P140 U1 ( .A1( _a[1] ), .A2( _a[9] ), .Z( _aa[1] ) );
XOR2UD1BWP30P140 U2 ( .A1( _a[2] ), .A2( _a[10] ), .Z( _aa[2] ) );
XOR2UD1BWP30P140 U3 ( .A1( _a[3] ), .A2( _a[11] ), .Z( _aa[3] ) );
XOR2UD1BWP30P140 U4 ( .A1( _a[4] ), .A2( _a[12] ), .Z( _aa[4] ) );
XOR2UD1BWP30P140 U5 ( .A1( _a[5] ), .A2( _a[13] ), .Z( _aa[5] ) );
XOR2UD1BWP30P140 U6 ( .A1( _a[6] ), .A2( _a[14] ), .Z( _aa[6] ) );
XOR2UD1BWP30P140 U7 ( .A1( _a[7] ), .A2( _a[15] ), .Z( _aa[7] ) );
XOR2UD1BWP30P140 U8 ( .A1( _b[0] ), .A2( _b[8] ), .Z( _bb[0] ) );
XOR2UD1BWP30P140 U9 ( .A1( _b[1] ), .A2( _b[9] ), .Z( _bb[1] ) );
XOR2UD1BWP30P140 U10 ( .A1( _b[2] ), .A2( _b[10] ), .Z( _bb[2] ) );
XOR2UD1BWP30P140 U11 ( .A1( _b[3] ), .A2( _b[11] ), .Z( _bb[3] ) );
XOR2UD1BWP30P140 U12 ( .A1( _b[4] ), .A2( _b[12] ), .Z( _bb[4] ) );
XOR2UD1BWP30P140 U13 ( .A1( _b[5] ), .A2( _b[13] ), .Z( _bb[5] ) );
XOR2UD1BWP30P140 U14 ( .A1( _b[6] ), .A2( _b[14] ), .Z( _bb[6] ) );
XOR2UD1BWP30P140 U15 ( .A1( _b[7] ), .A2( _b[15] ), .Z( _bb[7] ) );
endmodule
