module s_64bit ( a, b, aa, bb );
input [63:0] a;
input [63:0] b;
output [31:0] aa;
output [31:0] bb;
wire [31:0] _aa;
wire [31:0] _bb;
wire [63:0] _a;
wire [63:0] _b;
assign _a = a;
assign _b = b;
assign aa = _aa;
assign bb = _bb;
XOR2UD1BWP30P140 U0 ( .A1( _a[0] ), .A2( _a[32] ), .Z( _aa[0] ) );
XOR2UD1BWP30P140 U1 ( .A1( _a[1] ), .A2( _a[33] ), .Z( _aa[1] ) );
XOR2UD1BWP30P140 U2 ( .A1( _a[2] ), .A2( _a[34] ), .Z( _aa[2] ) );
XOR2UD1BWP30P140 U3 ( .A1( _a[3] ), .A2( _a[35] ), .Z( _aa[3] ) );
XOR2UD1BWP30P140 U4 ( .A1( _a[4] ), .A2( _a[36] ), .Z( _aa[4] ) );
XOR2UD1BWP30P140 U5 ( .A1( _a[5] ), .A2( _a[37] ), .Z( _aa[5] ) );
XOR2UD1BWP30P140 U6 ( .A1( _a[6] ), .A2( _a[38] ), .Z( _aa[6] ) );
XOR2UD1BWP30P140 U7 ( .A1( _a[7] ), .A2( _a[39] ), .Z( _aa[7] ) );
XOR2UD1BWP30P140 U8 ( .A1( _a[8] ), .A2( _a[40] ), .Z( _aa[8] ) );
XOR2UD1BWP30P140 U9 ( .A1( _a[9] ), .A2( _a[41] ), .Z( _aa[9] ) );
XOR2UD1BWP30P140 U10 ( .A1( _a[10] ), .A2( _a[42] ), .Z( _aa[10] ) );
XOR2UD1BWP30P140 U11 ( .A1( _a[11] ), .A2( _a[43] ), .Z( _aa[11] ) );
XOR2UD1BWP30P140 U12 ( .A1( _a[12] ), .A2( _a[44] ), .Z( _aa[12] ) );
XOR2UD1BWP30P140 U13 ( .A1( _a[13] ), .A2( _a[45] ), .Z( _aa[13] ) );
XOR2UD1BWP30P140 U14 ( .A1( _a[14] ), .A2( _a[46] ), .Z( _aa[14] ) );
XOR2UD1BWP30P140 U15 ( .A1( _a[15] ), .A2( _a[47] ), .Z( _aa[15] ) );
XOR2UD1BWP30P140 U16 ( .A1( _a[16] ), .A2( _a[48] ), .Z( _aa[16] ) );
XOR2UD1BWP30P140 U17 ( .A1( _a[17] ), .A2( _a[49] ), .Z( _aa[17] ) );
XOR2UD1BWP30P140 U18 ( .A1( _a[18] ), .A2( _a[50] ), .Z( _aa[18] ) );
XOR2UD1BWP30P140 U19 ( .A1( _a[19] ), .A2( _a[51] ), .Z( _aa[19] ) );
XOR2UD1BWP30P140 U20 ( .A1( _a[20] ), .A2( _a[52] ), .Z( _aa[20] ) );
XOR2UD1BWP30P140 U21 ( .A1( _a[21] ), .A2( _a[53] ), .Z( _aa[21] ) );
XOR2UD1BWP30P140 U22 ( .A1( _a[22] ), .A2( _a[54] ), .Z( _aa[22] ) );
XOR2UD1BWP30P140 U23 ( .A1( _a[23] ), .A2( _a[55] ), .Z( _aa[23] ) );
XOR2UD1BWP30P140 U24 ( .A1( _a[24] ), .A2( _a[56] ), .Z( _aa[24] ) );
XOR2UD1BWP30P140 U25 ( .A1( _a[25] ), .A2( _a[57] ), .Z( _aa[25] ) );
XOR2UD1BWP30P140 U26 ( .A1( _a[26] ), .A2( _a[58] ), .Z( _aa[26] ) );
XOR2UD1BWP30P140 U27 ( .A1( _a[27] ), .A2( _a[59] ), .Z( _aa[27] ) );
XOR2UD1BWP30P140 U28 ( .A1( _a[28] ), .A2( _a[60] ), .Z( _aa[28] ) );
XOR2UD1BWP30P140 U29 ( .A1( _a[29] ), .A2( _a[61] ), .Z( _aa[29] ) );
XOR2UD1BWP30P140 U30 ( .A1( _a[30] ), .A2( _a[62] ), .Z( _aa[30] ) );
XOR2UD1BWP30P140 U31 ( .A1( _a[31] ), .A2( _a[63] ), .Z( _aa[31] ) );
XOR2UD1BWP30P140 U32 ( .A1( _b[0] ), .A2( _b[32] ), .Z( _bb[0] ) );
XOR2UD1BWP30P140 U33 ( .A1( _b[1] ), .A2( _b[33] ), .Z( _bb[1] ) );
XOR2UD1BWP30P140 U34 ( .A1( _b[2] ), .A2( _b[34] ), .Z( _bb[2] ) );
XOR2UD1BWP30P140 U35 ( .A1( _b[3] ), .A2( _b[35] ), .Z( _bb[3] ) );
XOR2UD1BWP30P140 U36 ( .A1( _b[4] ), .A2( _b[36] ), .Z( _bb[4] ) );
XOR2UD1BWP30P140 U37 ( .A1( _b[5] ), .A2( _b[37] ), .Z( _bb[5] ) );
XOR2UD1BWP30P140 U38 ( .A1( _b[6] ), .A2( _b[38] ), .Z( _bb[6] ) );
XOR2UD1BWP30P140 U39 ( .A1( _b[7] ), .A2( _b[39] ), .Z( _bb[7] ) );
XOR2UD1BWP30P140 U40 ( .A1( _b[8] ), .A2( _b[40] ), .Z( _bb[8] ) );
XOR2UD1BWP30P140 U41 ( .A1( _b[9] ), .A2( _b[41] ), .Z( _bb[9] ) );
XOR2UD1BWP30P140 U42 ( .A1( _b[10] ), .A2( _b[42] ), .Z( _bb[10] ) );
XOR2UD1BWP30P140 U43 ( .A1( _b[11] ), .A2( _b[43] ), .Z( _bb[11] ) );
XOR2UD1BWP30P140 U44 ( .A1( _b[12] ), .A2( _b[44] ), .Z( _bb[12] ) );
XOR2UD1BWP30P140 U45 ( .A1( _b[13] ), .A2( _b[45] ), .Z( _bb[13] ) );
XOR2UD1BWP30P140 U46 ( .A1( _b[14] ), .A2( _b[46] ), .Z( _bb[14] ) );
XOR2UD1BWP30P140 U47 ( .A1( _b[15] ), .A2( _b[47] ), .Z( _bb[15] ) );
XOR2UD1BWP30P140 U48 ( .A1( _b[16] ), .A2( _b[48] ), .Z( _bb[16] ) );
XOR2UD1BWP30P140 U49 ( .A1( _b[17] ), .A2( _b[49] ), .Z( _bb[17] ) );
XOR2UD1BWP30P140 U50 ( .A1( _b[18] ), .A2( _b[50] ), .Z( _bb[18] ) );
XOR2UD1BWP30P140 U51 ( .A1( _b[19] ), .A2( _b[51] ), .Z( _bb[19] ) );
XOR2UD1BWP30P140 U52 ( .A1( _b[20] ), .A2( _b[52] ), .Z( _bb[20] ) );
XOR2UD1BWP30P140 U53 ( .A1( _b[21] ), .A2( _b[53] ), .Z( _bb[21] ) );
XOR2UD1BWP30P140 U54 ( .A1( _b[22] ), .A2( _b[54] ), .Z( _bb[22] ) );
XOR2UD1BWP30P140 U55 ( .A1( _b[23] ), .A2( _b[55] ), .Z( _bb[23] ) );
XOR2UD1BWP30P140 U56 ( .A1( _b[24] ), .A2( _b[56] ), .Z( _bb[24] ) );
XOR2UD1BWP30P140 U57 ( .A1( _b[25] ), .A2( _b[57] ), .Z( _bb[25] ) );
XOR2UD1BWP30P140 U58 ( .A1( _b[26] ), .A2( _b[58] ), .Z( _bb[26] ) );
XOR2UD1BWP30P140 U59 ( .A1( _b[27] ), .A2( _b[59] ), .Z( _bb[27] ) );
XOR2UD1BWP30P140 U60 ( .A1( _b[28] ), .A2( _b[60] ), .Z( _bb[28] ) );
XOR2UD1BWP30P140 U61 ( .A1( _b[29] ), .A2( _b[61] ), .Z( _bb[29] ) );
XOR2UD1BWP30P140 U62 ( .A1( _b[30] ), .A2( _b[62] ), .Z( _bb[30] ) );
XOR2UD1BWP30P140 U63 ( .A1( _b[31] ), .A2( _b[63] ), .Z( _bb[31] ) );
endmodule
