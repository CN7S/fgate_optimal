module gf_mul_128 ( a, b, c );
input [127:0] a;
input [127:0] b;
output [127:0] c;
wire [127:0] _c;
wire [127:0] _a;
wire [127:0] _b;
wire [254:0] d;
assign _a = a;
assign _b = b;
assign c = _c;
OKA_128bit mul_128_x ( .a( { _a[0], _a[1], _a[2], _a[3], _a[4], _a[5], _a[6], _a[7], _a[8], _a[9], _a[10], _a[11], _a[12], _a[13], _a[14], _a[15], _a[16], _a[17], _a[18], _a[19], _a[20], _a[21], _a[22], _a[23], _a[24], _a[25], _a[26], _a[27], _a[28], _a[29], _a[30], _a[31], _a[32], _a[33], _a[34], _a[35], _a[36], _a[37], _a[38], _a[39], _a[40], _a[41], _a[42], _a[43], _a[44], _a[45], _a[46], _a[47], _a[48], _a[49], _a[50], _a[51], _a[52], _a[53], _a[54], _a[55], _a[56], _a[57], _a[58], _a[59], _a[60], _a[61], _a[62], _a[63], _a[64], _a[65], _a[66], _a[67], _a[68], _a[69], _a[70], _a[71], _a[72], _a[73], _a[74], _a[75], _a[76], _a[77], _a[78], _a[79], _a[80], _a[81], _a[82], _a[83], _a[84], _a[85], _a[86], _a[87], _a[88], _a[89], _a[90], _a[91], _a[92], _a[93], _a[94], _a[95], _a[96], _a[97], _a[98], _a[99], _a[100], _a[101], _a[102], _a[103], _a[104], _a[105], _a[106], _a[107], _a[108], _a[109], _a[110], _a[111], _a[112], _a[113], _a[114], _a[115], _a[116], _a[117], _a[118], _a[119], _a[120], _a[121], _a[122], _a[123], _a[124], _a[125], _a[126], _a[127] } ), .b( { _b[0], _b[1], _b[2], _b[3], _b[4], _b[5], _b[6], _b[7], _b[8], _b[9], _b[10], _b[11], _b[12], _b[13], _b[14], _b[15], _b[16], _b[17], _b[18], _b[19], _b[20], _b[21], _b[22], _b[23], _b[24], _b[25], _b[26], _b[27], _b[28], _b[29], _b[30], _b[31], _b[32], _b[33], _b[34], _b[35], _b[36], _b[37], _b[38], _b[39], _b[40], _b[41], _b[42], _b[43], _b[44], _b[45], _b[46], _b[47], _b[48], _b[49], _b[50], _b[51], _b[52], _b[53], _b[54], _b[55], _b[56], _b[57], _b[58], _b[59], _b[60], _b[61], _b[62], _b[63], _b[64], _b[65], _b[66], _b[67], _b[68], _b[69], _b[70], _b[71], _b[72], _b[73], _b[74], _b[75], _b[76], _b[77], _b[78], _b[79], _b[80], _b[81], _b[82], _b[83], _b[84], _b[85], _b[86], _b[87], _b[88], _b[89], _b[90], _b[91], _b[92], _b[93], _b[94], _b[95], _b[96], _b[97], _b[98], _b[99], _b[100], _b[101], _b[102], _b[103], _b[104], _b[105], _b[106], _b[107], _b[108], _b[109], _b[110], _b[111], _b[112], _b[113], _b[114], _b[115], _b[116], _b[117], _b[118], _b[119], _b[120], _b[121], _b[122], _b[123], _b[124], _b[125], _b[126], _b[127] } ), .y( d ) );
reduction reduction_x ( .a( d ), .b( { _c[0], _c[1], _c[2], _c[3], _c[4], _c[5], _c[6], _c[7], _c[8], _c[9], _c[10], _c[11], _c[12], _c[13], _c[14], _c[15], _c[16], _c[17], _c[18], _c[19], _c[20], _c[21], _c[22], _c[23], _c[24], _c[25], _c[26], _c[27], _c[28], _c[29], _c[30], _c[31], _c[32], _c[33], _c[34], _c[35], _c[36], _c[37], _c[38], _c[39], _c[40], _c[41], _c[42], _c[43], _c[44], _c[45], _c[46], _c[47], _c[48], _c[49], _c[50], _c[51], _c[52], _c[53], _c[54], _c[55], _c[56], _c[57], _c[58], _c[59], _c[60], _c[61], _c[62], _c[63], _c[64], _c[65], _c[66], _c[67], _c[68], _c[69], _c[70], _c[71], _c[72], _c[73], _c[74], _c[75], _c[76], _c[77], _c[78], _c[79], _c[80], _c[81], _c[82], _c[83], _c[84], _c[85], _c[86], _c[87], _c[88], _c[89], _c[90], _c[91], _c[92], _c[93], _c[94], _c[95], _c[96], _c[97], _c[98], _c[99], _c[100], _c[101], _c[102], _c[103], _c[104], _c[105], _c[106], _c[107], _c[108], _c[109], _c[110], _c[111], _c[112], _c[113], _c[114], _c[115], _c[116], _c[117], _c[118], _c[119], _c[120], _c[121], _c[122], _c[123], _c[124], _c[125], _c[126], _c[127] } ) );
endmodule
