module OKA_128bit ( a, b, y, C_g1, rst_n );
input [127:0] a;
input [127:0] b;
output [254:0] y;
input [21:0] C_g1;
input rst_n;
wire [254:0] _y;
wire [21:0] _C_g1;
wire [63:0] aa;
wire [63:0] bb;
wire [63:0] al;
wire [63:0] ah;
wire [63:0] bl;
wire [63:0] bh;
wire [126:0] z0;
wire [126:0] z1;
wire [126:0] z2;
wire _rst_n;
assign al[0] = a[0];
assign ah[0] = a[1];
assign al[1] = a[2];
assign ah[1] = a[3];
assign al[2] = a[4];
assign ah[2] = a[5];
assign al[3] = a[6];
assign ah[3] = a[7];
assign al[4] = a[8];
assign ah[4] = a[9];
assign al[5] = a[10];
assign ah[5] = a[11];
assign al[6] = a[12];
assign ah[6] = a[13];
assign al[7] = a[14];
assign ah[7] = a[15];
assign al[8] = a[16];
assign ah[8] = a[17];
assign al[9] = a[18];
assign ah[9] = a[19];
assign al[10] = a[20];
assign ah[10] = a[21];
assign al[11] = a[22];
assign ah[11] = a[23];
assign al[12] = a[24];
assign ah[12] = a[25];
assign al[13] = a[26];
assign ah[13] = a[27];
assign al[14] = a[28];
assign ah[14] = a[29];
assign al[15] = a[30];
assign ah[15] = a[31];
assign al[16] = a[32];
assign ah[16] = a[33];
assign al[17] = a[34];
assign ah[17] = a[35];
assign al[18] = a[36];
assign ah[18] = a[37];
assign al[19] = a[38];
assign ah[19] = a[39];
assign al[20] = a[40];
assign ah[20] = a[41];
assign al[21] = a[42];
assign ah[21] = a[43];
assign al[22] = a[44];
assign ah[22] = a[45];
assign al[23] = a[46];
assign ah[23] = a[47];
assign al[24] = a[48];
assign ah[24] = a[49];
assign al[25] = a[50];
assign ah[25] = a[51];
assign al[26] = a[52];
assign ah[26] = a[53];
assign al[27] = a[54];
assign ah[27] = a[55];
assign al[28] = a[56];
assign ah[28] = a[57];
assign al[29] = a[58];
assign ah[29] = a[59];
assign al[30] = a[60];
assign ah[30] = a[61];
assign al[31] = a[62];
assign ah[31] = a[63];
assign al[32] = a[64];
assign ah[32] = a[65];
assign al[33] = a[66];
assign ah[33] = a[67];
assign al[34] = a[68];
assign ah[34] = a[69];
assign al[35] = a[70];
assign ah[35] = a[71];
assign al[36] = a[72];
assign ah[36] = a[73];
assign al[37] = a[74];
assign ah[37] = a[75];
assign al[38] = a[76];
assign ah[38] = a[77];
assign al[39] = a[78];
assign ah[39] = a[79];
assign al[40] = a[80];
assign ah[40] = a[81];
assign al[41] = a[82];
assign ah[41] = a[83];
assign al[42] = a[84];
assign ah[42] = a[85];
assign al[43] = a[86];
assign ah[43] = a[87];
assign al[44] = a[88];
assign ah[44] = a[89];
assign al[45] = a[90];
assign ah[45] = a[91];
assign al[46] = a[92];
assign ah[46] = a[93];
assign al[47] = a[94];
assign ah[47] = a[95];
assign al[48] = a[96];
assign ah[48] = a[97];
assign al[49] = a[98];
assign ah[49] = a[99];
assign al[50] = a[100];
assign ah[50] = a[101];
assign al[51] = a[102];
assign ah[51] = a[103];
assign al[52] = a[104];
assign ah[52] = a[105];
assign al[53] = a[106];
assign ah[53] = a[107];
assign al[54] = a[108];
assign ah[54] = a[109];
assign al[55] = a[110];
assign ah[55] = a[111];
assign al[56] = a[112];
assign ah[56] = a[113];
assign al[57] = a[114];
assign ah[57] = a[115];
assign al[58] = a[116];
assign ah[58] = a[117];
assign al[59] = a[118];
assign ah[59] = a[119];
assign al[60] = a[120];
assign ah[60] = a[121];
assign al[61] = a[122];
assign ah[61] = a[123];
assign al[62] = a[124];
assign ah[62] = a[125];
assign al[63] = a[126];
assign ah[63] = a[127];
assign bl[0] = b[0];
assign bh[0] = b[1];
assign bl[1] = b[2];
assign bh[1] = b[3];
assign bl[2] = b[4];
assign bh[2] = b[5];
assign bl[3] = b[6];
assign bh[3] = b[7];
assign bl[4] = b[8];
assign bh[4] = b[9];
assign bl[5] = b[10];
assign bh[5] = b[11];
assign bl[6] = b[12];
assign bh[6] = b[13];
assign bl[7] = b[14];
assign bh[7] = b[15];
assign bl[8] = b[16];
assign bh[8] = b[17];
assign bl[9] = b[18];
assign bh[9] = b[19];
assign bl[10] = b[20];
assign bh[10] = b[21];
assign bl[11] = b[22];
assign bh[11] = b[23];
assign bl[12] = b[24];
assign bh[12] = b[25];
assign bl[13] = b[26];
assign bh[13] = b[27];
assign bl[14] = b[28];
assign bh[14] = b[29];
assign bl[15] = b[30];
assign bh[15] = b[31];
assign bl[16] = b[32];
assign bh[16] = b[33];
assign bl[17] = b[34];
assign bh[17] = b[35];
assign bl[18] = b[36];
assign bh[18] = b[37];
assign bl[19] = b[38];
assign bh[19] = b[39];
assign bl[20] = b[40];
assign bh[20] = b[41];
assign bl[21] = b[42];
assign bh[21] = b[43];
assign bl[22] = b[44];
assign bh[22] = b[45];
assign bl[23] = b[46];
assign bh[23] = b[47];
assign bl[24] = b[48];
assign bh[24] = b[49];
assign bl[25] = b[50];
assign bh[25] = b[51];
assign bl[26] = b[52];
assign bh[26] = b[53];
assign bl[27] = b[54];
assign bh[27] = b[55];
assign bl[28] = b[56];
assign bh[28] = b[57];
assign bl[29] = b[58];
assign bh[29] = b[59];
assign bl[30] = b[60];
assign bh[30] = b[61];
assign bl[31] = b[62];
assign bh[31] = b[63];
assign bl[32] = b[64];
assign bh[32] = b[65];
assign bl[33] = b[66];
assign bh[33] = b[67];
assign bl[34] = b[68];
assign bh[34] = b[69];
assign bl[35] = b[70];
assign bh[35] = b[71];
assign bl[36] = b[72];
assign bh[36] = b[73];
assign bl[37] = b[74];
assign bh[37] = b[75];
assign bl[38] = b[76];
assign bh[38] = b[77];
assign bl[39] = b[78];
assign bh[39] = b[79];
assign bl[40] = b[80];
assign bh[40] = b[81];
assign bl[41] = b[82];
assign bh[41] = b[83];
assign bl[42] = b[84];
assign bh[42] = b[85];
assign bl[43] = b[86];
assign bh[43] = b[87];
assign bl[44] = b[88];
assign bh[44] = b[89];
assign bl[45] = b[90];
assign bh[45] = b[91];
assign bl[46] = b[92];
assign bh[46] = b[93];
assign bl[47] = b[94];
assign bh[47] = b[95];
assign bl[48] = b[96];
assign bh[48] = b[97];
assign bl[49] = b[98];
assign bh[49] = b[99];
assign bl[50] = b[100];
assign bh[50] = b[101];
assign bl[51] = b[102];
assign bh[51] = b[103];
assign bl[52] = b[104];
assign bh[52] = b[105];
assign bl[53] = b[106];
assign bh[53] = b[107];
assign bl[54] = b[108];
assign bh[54] = b[109];
assign bl[55] = b[110];
assign bh[55] = b[111];
assign bl[56] = b[112];
assign bh[56] = b[113];
assign bl[57] = b[114];
assign bh[57] = b[115];
assign bl[58] = b[116];
assign bh[58] = b[117];
assign bl[59] = b[118];
assign bh[59] = b[119];
assign bl[60] = b[120];
assign bh[60] = b[121];
assign bl[61] = b[122];
assign bh[61] = b[123];
assign bl[62] = b[124];
assign bh[62] = b[125];
assign bl[63] = b[126];
assign bh[63] = b[127];
assign y = _y;
assign _C_g1 = C_g1;
assign _rst_n = rst_n;
s_128bit s128_u ( .a( { ah[63], al[63], ah[62], al[62], ah[61], al[61], ah[60], al[60], ah[59], al[59], ah[58], al[58], ah[57], al[57], ah[56], al[56], ah[55], al[55], ah[54], al[54], ah[53], al[53], ah[52], al[52], ah[51], al[51], ah[50], al[50], ah[49], al[49], ah[48], al[48], ah[47], al[47], ah[46], al[46], ah[45], al[45], ah[44], al[44], ah[43], al[43], ah[42], al[42], ah[41], al[41], ah[40], al[40], ah[39], al[39], ah[38], al[38], ah[37], al[37], ah[36], al[36], ah[35], al[35], ah[34], al[34], ah[33], al[33], ah[32], al[32], ah[31], al[31], ah[30], al[30], ah[29], al[29], ah[28], al[28], ah[27], al[27], ah[26], al[26], ah[25], al[25], ah[24], al[24], ah[23], al[23], ah[22], al[22], ah[21], al[21], ah[20], al[20], ah[19], al[19], ah[18], al[18], ah[17], al[17], ah[16], al[16], ah[15], al[15], ah[14], al[14], ah[13], al[13], ah[12], al[12], ah[11], al[11], ah[10], al[10], ah[9], al[9], ah[8], al[8], ah[7], al[7], ah[6], al[6], ah[5], al[5], ah[4], al[4], ah[3], al[3], ah[2], al[2], ah[1], al[1], ah[0], al[0] } ), .b( { bh[63], bl[63], bh[62], bl[62], bh[61], bl[61], bh[60], bl[60], bh[59], bl[59], bh[58], bl[58], bh[57], bl[57], bh[56], bl[56], bh[55], bl[55], bh[54], bl[54], bh[53], bl[53], bh[52], bl[52], bh[51], bl[51], bh[50], bl[50], bh[49], bl[49], bh[48], bl[48], bh[47], bl[47], bh[46], bl[46], bh[45], bl[45], bh[44], bl[44], bh[43], bl[43], bh[42], bl[42], bh[41], bl[41], bh[40], bl[40], bh[39], bl[39], bh[38], bl[38], bh[37], bl[37], bh[36], bl[36], bh[35], bl[35], bh[34], bl[34], bh[33], bl[33], bh[32], bl[32], bh[31], bl[31], bh[30], bl[30], bh[29], bl[29], bh[28], bl[28], bh[27], bl[27], bh[26], bl[26], bh[25], bl[25], bh[24], bl[24], bh[23], bl[23], bh[22], bl[22], bh[21], bl[21], bh[20], bl[20], bh[19], bl[19], bh[18], bl[18], bh[17], bl[17], bh[16], bl[16], bh[15], bl[15], bh[14], bl[14], bh[13], bl[13], bh[12], bl[12], bh[11], bl[11], bh[10], bl[10], bh[9], bl[9], bh[8], bl[8], bh[7], bl[7], bh[6], bl[6], bh[5], bl[5], bh[4], bl[4], bh[3], bl[3], bh[2], bl[2], bh[1], bl[1], bh[0], bl[0] } ), .aa( aa ), .bb( bb ) );
OKA_64bit mul64_0 ( .a( al ), .b( bl ), .y( z0 ), .C_g1( _C_g1 ), .rst_n( _rst_n ) );
OKA_64bit mul64_1 ( .a( aa ), .b( bb ), .y( z1 ), .C_g1( _C_g1 ), .rst_n( _rst_n ) );
OKA_64bit mul64_2 ( .a( ah ), .b( bh ), .y( z2 ), .C_g1( _C_g1 ), .rst_n( _rst_n ) );
os_128bit os128_u ( .z0( z0 ), .z1( z1 ), .z2( z2 ), .y( _y ), .C_g1( _C_g1 ), .rst_n( _rst_n ) );
endmodule
