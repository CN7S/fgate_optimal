module FXOR2UD1BWP30P140 (
    A1,A2,Z,en
);
    input A1;
    input A2;
    input en;
    output Z;
endmodule

module FXOR3UD1BWP30P140 (
    A1,A2,A3,Z,en
);
    input A1;
    input A2;
    input A3;
    input en;
    output Z;
endmodule
module FXOR4D1BWP30P140 (
    A1,A2,A3,A4,Z,en
);
    input A1;
    input A2;
    input A3;
    input A4;
    input en;
    output Z;
endmodule

module FCKND2D1BWP30P140 (
    A1,A2,ZN,en
);
    input A1;
    input A2;
    input en;
    output ZN;
endmodule

module FNR2D1BWP30P140 (
    A1,A2,ZN,en
);
    input A1;
    input A2;
    input en;
    output ZN;
endmodule
module FAN2D1BWP30P140 (
    A1,A2,Z,en
);
    input A1;
    input A2;
    input en;
    output Z;
endmodule
module FINR2D1BWP30P140 (
    A1,B1,ZN,en
);
    input A1;
    input B1;
    input en;
    output ZN;
endmodule
module FINVD1BWP30P140 (
    I,ZN,en
);
    input I;
    input en;
    output ZN;
endmodule
module FXNR3UD1BWP30P140 (
    A1,A2,A3,ZN,en
);
    input A1,A2,A3;
    input en;
    output ZN;
endmodule

module FXNR2UD1BWP30P140 (
    A1,A2,ZN,en
);
    input A1,A2;
    input en;
    output ZN;
endmodule