module reduction ( a, b, C_g1, rst_n );
  input [254:0] a;
  input [21:0] C_g1;
  input rst_n;
  output [127:0] b;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, b_98_, n14, b_96_,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, b_68_,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, b_45_, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, b_20_, n50, b_18_, n52, n53, b_14_,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145;
  assign b[98] = b_98_;
  assign b[96] = b_96_;
  assign b[68] = b_68_;
  assign b[45] = b_45_;
  assign b[20] = b_20_;
  assign b[18] = b_18_;
  assign b[14] = b_14_;

  XOR2UD1BWP30P140 U1 ( .A1(a[252]), .A2(a[131]), .Z(n97) );
  XOR2UD1BWP30P140 U2 ( .A1(a[253]), .A2(a[254]), .Z(n98) );
  XOR2UD1BWP30P140 U3 ( .A1(a[132]), .A2(a[253]), .Z(n104) );
  XOR2UD1BWP30P140 U4 ( .A1(a[129]), .A2(a[250]), .Z(n76) );
  XOR2UD1BWP30P140 U5 ( .A1(n6), .A2(a[240]), .Z(n139) );
  XNR2UD1BWP30P140 U6 ( .A1(a[250]), .A2(a[251]), .ZN(n118) );
  XOR2UD1BWP30P140 U7 ( .A1(n7), .A2(a[238]), .Z(n140) );
  XOR2UD1BWP30P140 U8 ( .A1(n8), .A2(a[236]), .Z(n141) );
  XOR2UD1BWP30P140 U9 ( .A1(n9), .A2(a[234]), .Z(n142) );
  XOR2UD1BWP30P140 U10 ( .A1(n10), .A2(a[232]), .Z(n143) );
  XOR2UD1BWP30P140 U11 ( .A1(n11), .A2(a[230]), .Z(n144) );
  XOR2UD1BWP30P140 U12 ( .A1(n12), .A2(a[228]), .Z(n145) );
  XOR2UD1BWP30P140 U13 ( .A1(n14), .A2(a[226]), .Z(n69) );
  XNR2UD1BWP30P140 U14 ( .A1(a[163]), .A2(a[164]), .ZN(n113) );
  XOR2UD1BWP30P140 U15 ( .A1(a[133]), .A2(a[134]), .Z(n82) );
  XOR2UD1BWP30P140 U16 ( .A1(a[135]), .A2(a[136]), .Z(n67) );
  XOR2UD1BWP30P140 U17 ( .A1(a[139]), .A2(a[140]), .Z(n130) );
  XNR2UD1BWP30P140 U18 ( .A1(a[186]), .A2(a[187]), .ZN(n96) );
  XOR2UD1BWP30P140 U19 ( .A1(n16), .A2(a[224]), .Z(n71) );
  XNR2UD1BWP30P140 U20 ( .A1(a[241]), .A2(a[242]), .ZN(n138) );
  XOR2UD1BWP30P140 U21 ( .A1(n19), .A2(a[214]), .Z(n78) );
  XOR2UD1BWP30P140 U22 ( .A1(n22), .A2(a[208]), .Z(n81) );
  XOR2UD1BWP30P140 U23 ( .A1(n29), .A2(a[196]), .Z(n90) );
  XOR2UD1BWP30P140 U24 ( .A1(n30), .A2(a[194]), .Z(n92) );
  XOR2UD1BWP30P140 U25 ( .A1(n23), .A2(a[206]), .Z(n84) );
  XOR2UD1BWP30P140 U26 ( .A1(n24), .A2(a[204]), .Z(n85) );
  XOR2UD1BWP30P140 U27 ( .A1(n25), .A2(a[202]), .Z(n86) );
  XOR2UD1BWP30P140 U28 ( .A1(n26), .A2(a[200]), .Z(n87) );
  XOR2UD1BWP30P140 U29 ( .A1(n27), .A2(a[198]), .Z(n88) );
  XOR2UD1BWP30P140 U30 ( .A1(n18), .A2(a[216]), .Z(n77) );
  XOR2UD1BWP30P140 U31 ( .A1(n20), .A2(a[212]), .Z(n79) );
  XOR2UD1BWP30P140 U32 ( .A1(n21), .A2(a[210]), .Z(n80) );
  XNR2UD1BWP30P140 U33 ( .A1(n83), .A2(a[254]), .ZN(n117) );
  XOR2UD1BWP30P140 U34 ( .A1(n17), .A2(a[222]), .Z(n73) );
  XOR2UD1BWP30P140 U35 ( .A1(n31), .A2(a[192]), .Z(n93) );
  XOR2UD1BWP30P140 U36 ( .A1(n43), .A2(a[160]), .Z(n115) );
  XOR2UD1BWP30P140 U37 ( .A1(n44), .A2(a[158]), .Z(n116) );
  XOR2UD1BWP30P140 U38 ( .A1(n45), .A2(a[156]), .Z(n119) );
  XOR2UD1BWP30P140 U39 ( .A1(n46), .A2(a[154]), .Z(n120) );
  XOR2UD1BWP30P140 U40 ( .A1(n47), .A2(a[152]), .Z(n121) );
  XOR2UD1BWP30P140 U41 ( .A1(n48), .A2(a[150]), .Z(n122) );
  XOR2UD1BWP30P140 U42 ( .A1(n50), .A2(a[148]), .Z(n123) );
  XOR2UD1BWP30P140 U43 ( .A1(n52), .A2(a[146]), .Z(n125) );
  XOR2UD1BWP30P140 U44 ( .A1(n53), .A2(a[144]), .Z(n127) );
  XNR2UD1BWP30P140 U45 ( .A1(a[219]), .A2(a[220]), .ZN(n74) );
  XNR2UD1BWP30P140 U46 ( .A1(a[217]), .A2(a[218]), .ZN(n75) );
  XOR2UD1BWP30P140 U47 ( .A1(a[130]), .A2(a[251]), .Z(n68) );
  XNR2UD1BWP30P140 U48 ( .A1(a[243]), .A2(a[244]), .ZN(n137) );
  XNR2UD1BWP30P140 U49 ( .A1(a[161]), .A2(a[162]), .ZN(n114) );
  XNR2UD1BWP30P140 U50 ( .A1(a[141]), .A2(a[142]), .ZN(n128) );
  XNR2UD1BWP30P140 U51 ( .A1(a[189]), .A2(a[190]), .ZN(n94) );
  XOR2UD1BWP30P140 U52 ( .A1(n34), .A2(a[181]), .Z(n101) );
  XOR2UD1BWP30P140 U53 ( .A1(n37), .A2(a[175]), .Z(n105) );
  XOR2UD1BWP30P140 U54 ( .A1(n39), .A2(a[173]), .Z(n106) );
  XOR2UD1BWP30P140 U55 ( .A1(n40), .A2(a[171]), .Z(n108) );
  XOR2UD1BWP30P140 U56 ( .A1(n41), .A2(a[169]), .Z(n109) );
  XOR2UD1BWP30P140 U57 ( .A1(n33), .A2(a[183]), .Z(n100) );
  XOR2UD1BWP30P140 U58 ( .A1(n35), .A2(a[179]), .Z(n102) );
  XOR2UD1BWP30P140 U59 ( .A1(n36), .A2(a[177]), .Z(n103) );
  XNR2UD1BWP30P140 U60 ( .A1(a[246]), .A2(a[247]), .ZN(n134) );
  XNR2UD1BWP30P140 U61 ( .A1(n98), .A2(a[132]), .ZN(n89) );
  XOR2UD1BWP30P140 U62 ( .A1(a[137]), .A2(a[138]), .Z(n135) );
  XNR2UD1BWP30P140 U63 ( .A1(a[184]), .A2(a[185]), .ZN(n99) );
  XNR2UD1BWP30P140 U64 ( .A1(a[166]), .A2(a[167]), .ZN(n110) );
  XNR2UD1BWP30P140 U65 ( .A1(n1), .A2(a[128]), .ZN(n83) );
  XOR2UD1BWP30P140 U66 ( .A1(a[248]), .A2(n1), .Z(n133) );
  XNR2UD1BWP30P140 U67 ( .A1(a[0]), .A2(n117), .ZN(b[0]) );
  INVD1BWP30P140 U68 ( .I(a[245]), .ZN(n3) );
  INVD1BWP30P140 U69 ( .I(a[249]), .ZN(n1) );
  INVD1BWP30P140 U70 ( .I(a[239]), .ZN(n6) );
  INVD1BWP30P140 U71 ( .I(a[237]), .ZN(n7) );
  INVD1BWP30P140 U72 ( .I(a[235]), .ZN(n8) );
  INVD1BWP30P140 U73 ( .I(a[233]), .ZN(n9) );
  INVD1BWP30P140 U74 ( .I(a[231]), .ZN(n10) );
  INVD1BWP30P140 U75 ( .I(a[229]), .ZN(n11) );
  INVD1BWP30P140 U76 ( .I(n107), .ZN(b_45_) );
  XOR4D1BWP30P140 U77 ( .A1(a[45]), .A2(a[171]), .A3(a[166]), .A4(n106), .Z(
        n107) );
  INVD1BWP30P140 U78 ( .I(n91), .ZN(b_68_) );
  XOR4D1BWP30P140 U79 ( .A1(a[68]), .A2(a[194]), .A3(a[189]), .A4(n90), .Z(n91) );
  INVD1BWP30P140 U80 ( .I(n70), .ZN(b_98_) );
  XOR4D1BWP30P140 U81 ( .A1(a[98]), .A2(a[224]), .A3(a[219]), .A4(n69), .Z(n70) );
  INVD1BWP30P140 U82 ( .I(n72), .ZN(b_96_) );
  XOR4D1BWP30P140 U83 ( .A1(a[96]), .A2(a[222]), .A3(a[217]), .A4(n71), .Z(n72) );
  INVD1BWP30P140 U84 ( .I(a[182]), .ZN(n33) );
  XOR4D1BWP30P140 U85 ( .A1(a[252]), .A2(a[126]), .A3(a[247]), .A4(n98), .Z(
        b[126]) );
  XOR4D1BWP30P140 U86 ( .A1(a[252]), .A2(a[124]), .A3(n3), .A4(n118), .Z(
        b[124]) );
  INVD1BWP30P140 U87 ( .I(a[176]), .ZN(n36) );
  INVD1BWP30P140 U88 ( .I(a[174]), .ZN(n37) );
  INVD1BWP30P140 U89 ( .I(a[170]), .ZN(n40) );
  INVD1BWP30P140 U90 ( .I(a[168]), .ZN(n41) );
  INVD1BWP30P140 U91 ( .I(a[180]), .ZN(n34) );
  INVD1BWP30P140 U92 ( .I(a[178]), .ZN(n35) );
  INVD1BWP30P140 U93 ( .I(a[227]), .ZN(n12) );
  INVD1BWP30P140 U94 ( .I(a[225]), .ZN(n14) );
  INVD1BWP30P140 U95 ( .I(a[223]), .ZN(n16) );
  XOR4D1BWP30P140 U96 ( .A1(n65), .A2(a[142]), .A3(a[137]), .A4(n127), .Z(
        b[16]) );
  INVD1BWP30P140 U97 ( .I(a[16]), .ZN(n65) );
  XOR4D1BWP30P140 U98 ( .A1(n66), .A2(n97), .A3(a[133]), .A4(n89), .Z(b[5]) );
  INVD1BWP30P140 U99 ( .I(a[5]), .ZN(n66) );
  XOR4D1BWP30P140 U100 ( .A1(n63), .A2(a[163]), .A3(a[156]), .A4(n114), .Z(
        b[35]) );
  INVD1BWP30P140 U101 ( .I(a[35]), .ZN(n63) );
  XOR4D1BWP30P140 U102 ( .A1(n59), .A2(a[186]), .A3(a[179]), .A4(n99), .Z(
        b[58]) );
  INVD1BWP30P140 U103 ( .I(a[58]), .ZN(n59) );
  XOR4D1BWP30P140 U104 ( .A1(n60), .A2(a[184]), .A3(a[177]), .A4(n100), .Z(
        b[56]) );
  INVD1BWP30P140 U105 ( .I(a[56]), .ZN(n60) );
  XOR4D1BWP30P140 U106 ( .A1(n64), .A2(a[161]), .A3(a[154]), .A4(n115), .Z(
        b[33]) );
  INVD1BWP30P140 U107 ( .I(a[33]), .ZN(n64) );
  XOR4D1BWP30P140 U108 ( .A1(n61), .A2(a[169]), .A3(a[164]), .A4(n108), .Z(
        b[43]) );
  INVD1BWP30P140 U109 ( .I(a[43]), .ZN(n61) );
  XOR4D1BWP30P140 U110 ( .A1(n62), .A2(a[167]), .A3(a[162]), .A4(n109), .Z(
        b[41]) );
  INVD1BWP30P140 U111 ( .I(a[41]), .ZN(n62) );
  XOR4D1BWP30P140 U112 ( .A1(n58), .A2(a[190]), .A3(a[185]), .A4(n93), .Z(
        b[64]) );
  INVD1BWP30P140 U113 ( .I(a[64]), .ZN(n58) );
  XOR4D1BWP30P140 U114 ( .A1(n55), .A2(a[219]), .A3(a[212]), .A4(n75), .Z(
        b[91]) );
  INVD1BWP30P140 U115 ( .I(a[91]), .ZN(n55) );
  XOR4D1BWP30P140 U116 ( .A1(n56), .A2(a[217]), .A3(a[210]), .A4(n77), .Z(
        b[89]) );
  INVD1BWP30P140 U117 ( .I(a[89]), .ZN(n56) );
  XOR4D1BWP30P140 U118 ( .A1(n2), .A2(a[121]), .A3(a[242]), .A4(n133), .Z(
        b[121]) );
  INVD1BWP30P140 U119 ( .I(a[247]), .ZN(n2) );
  XOR4D1BWP30P140 U120 ( .A1(n57), .A2(a[192]), .A3(a[187]), .A4(n92), .Z(
        b[66]) );
  INVD1BWP30P140 U121 ( .I(a[66]), .ZN(n57) );
  XOR4D1BWP30P140 U122 ( .A1(n4), .A2(a[115]), .A3(a[236]), .A4(n138), .Z(
        b[115]) );
  XOR4D1BWP30P140 U123 ( .A1(n5), .A2(a[113]), .A3(a[234]), .A4(n139), .Z(
        b[113]) );
  XOR4D1BWP30P140 U124 ( .A1(n7), .A2(a[109]), .A3(a[230]), .A4(n141), .Z(
        b[109]) );
  XOR4D1BWP30P140 U125 ( .A1(n8), .A2(a[107]), .A3(a[228]), .A4(n142), .Z(
        b[107]) );
  XOR4D1BWP30P140 U126 ( .A1(n9), .A2(a[105]), .A3(a[226]), .A4(n143), .Z(
        b[105]) );
  XOR4D1BWP30P140 U127 ( .A1(n10), .A2(a[103]), .A3(a[224]), .A4(n144), .Z(
        b[103]) );
  XOR4D1BWP30P140 U128 ( .A1(n11), .A2(a[101]), .A3(a[222]), .A4(n145), .Z(
        b[101]) );
  XOR4D1BWP30P140 U129 ( .A1(n6), .A2(a[111]), .A3(a[232]), .A4(n140), .Z(
        b[111]) );
  XOR4D1BWP30P140 U130 ( .A1(n1), .A2(a[123]), .A3(a[244]), .A4(n118), .Z(
        b[123]) );
  XOR4D1BWP30P140 U131 ( .A1(n3), .A2(a[119]), .A3(a[240]), .A4(n134), .Z(
        b[119]) );
  XOR4D1BWP30P140 U132 ( .A1(n3), .A2(a[117]), .A3(a[238]), .A4(n137), .Z(
        b[117]) );
  XOR4D1BWP30P140 U133 ( .A1(n136), .A2(a[118]), .A3(a[244]), .A4(a[239]), .Z(
        b[118]) );
  XNR2UD1BWP30P140 U134 ( .A1(a[246]), .A2(n3), .ZN(n136) );
  XOR4D1BWP30P140 U135 ( .A1(a[250]), .A2(a[122]), .A3(n4), .A4(n133), .Z(
        b[122]) );
  XOR4D1BWP30P140 U136 ( .A1(n112), .A2(a[38]), .A3(a[166]), .A4(a[165]), .Z(
        b[38]) );
  XOR2UD1BWP30P140 U137 ( .A1(a[164]), .A2(a[159]), .Z(n112) );
  XOR4D1BWP30P140 U138 ( .A1(a[99]), .A2(n12), .A3(a[220]), .A4(n69), .Z(b[99]) );
  XOR4D1BWP30P140 U139 ( .A1(a[97]), .A2(n14), .A3(a[218]), .A4(n71), .Z(b[97]) );
  XOR4D1BWP30P140 U140 ( .A1(a[93]), .A2(n17), .A3(a[214]), .A4(n74), .Z(b[93]) );
  XOR4D1BWP30P140 U141 ( .A1(a[73]), .A2(n25), .A3(a[194]), .A4(n87), .Z(b[73]) );
  XOR4D1BWP30P140 U142 ( .A1(a[69]), .A2(n27), .A3(a[190]), .A4(n90), .Z(b[69]) );
  XOR4D1BWP30P140 U143 ( .A1(a[67]), .A2(a[195]), .A3(n32), .A4(n92), .Z(b[67]) );
  XOR4D1BWP30P140 U144 ( .A1(a[65]), .A2(n30), .A3(a[186]), .A4(n93), .Z(b[65]) );
  XOR4D1BWP30P140 U145 ( .A1(a[95]), .A2(n16), .A3(a[216]), .A4(n73), .Z(b[95]) );
  XOR4D1BWP30P140 U146 ( .A1(a[87]), .A2(n18), .A3(a[208]), .A4(n78), .Z(b[87]) );
  XOR4D1BWP30P140 U147 ( .A1(a[85]), .A2(n19), .A3(a[206]), .A4(n79), .Z(b[85]) );
  XOR4D1BWP30P140 U148 ( .A1(a[83]), .A2(n20), .A3(a[204]), .A4(n80), .Z(b[83]) );
  XOR4D1BWP30P140 U149 ( .A1(a[81]), .A2(n21), .A3(a[202]), .A4(n81), .Z(b[81]) );
  XOR4D1BWP30P140 U150 ( .A1(a[79]), .A2(n22), .A3(a[200]), .A4(n84), .Z(b[79]) );
  XOR4D1BWP30P140 U151 ( .A1(a[77]), .A2(n23), .A3(a[198]), .A4(n85), .Z(b[77]) );
  XOR4D1BWP30P140 U152 ( .A1(a[75]), .A2(n24), .A3(a[196]), .A4(n86), .Z(b[75]) );
  XOR4D1BWP30P140 U153 ( .A1(a[71]), .A2(n26), .A3(a[192]), .A4(n88), .Z(b[71]) );
  XOR4D1BWP30P140 U154 ( .A1(n95), .A2(a[61]), .A3(a[189]), .A4(a[188]), .Z(
        b[61]) );
  XOR2UD1BWP30P140 U155 ( .A1(a[187]), .A2(a[182]), .Z(n95) );
  XOR4D1BWP30P140 U156 ( .A1(a[63]), .A2(n31), .A3(a[184]), .A4(n94), .Z(b[63]) );
  XOR4D1BWP30P140 U157 ( .A1(a[59]), .A2(a[185]), .A3(n34), .A4(n96), .Z(b[59]) );
  XOR4D1BWP30P140 U158 ( .A1(a[57]), .A2(a[183]), .A3(n35), .A4(n99), .Z(b[57]) );
  XOR4D1BWP30P140 U159 ( .A1(a[55]), .A2(a[181]), .A3(n36), .A4(n100), .Z(
        b[55]) );
  XOR4D1BWP30P140 U160 ( .A1(a[53]), .A2(a[179]), .A3(n37), .A4(n101), .Z(
        b[53]) );
  XOR4D1BWP30P140 U161 ( .A1(a[37]), .A2(n42), .A3(a[158]), .A4(n113), .Z(
        b[37]) );
  XOR4D1BWP30P140 U162 ( .A1(a[51]), .A2(a[177]), .A3(n39), .A4(n102), .Z(
        b[51]) );
  XOR4D1BWP30P140 U163 ( .A1(a[49]), .A2(a[175]), .A3(n40), .A4(n103), .Z(
        b[49]) );
  XOR4D1BWP30P140 U164 ( .A1(a[47]), .A2(a[173]), .A3(n41), .A4(n105), .Z(
        b[47]) );
  XOR4D1BWP30P140 U165 ( .A1(a[39]), .A2(n42), .A3(a[160]), .A4(n110), .Z(
        b[39]) );
  INVD1BWP30P140 U166 ( .I(a[159]), .ZN(n43) );
  XOR4D1BWP30P140 U167 ( .A1(a[31]), .A2(n43), .A3(a[152]), .A4(n116), .Z(
        b[31]) );
  XOR4D1BWP30P140 U168 ( .A1(a[29]), .A2(n44), .A3(a[150]), .A4(n119), .Z(
        b[29]) );
  XOR4D1BWP30P140 U169 ( .A1(a[27]), .A2(n45), .A3(a[148]), .A4(n120), .Z(
        b[27]) );
  XOR4D1BWP30P140 U170 ( .A1(a[25]), .A2(n46), .A3(a[146]), .A4(n121), .Z(
        b[25]) );
  XOR4D1BWP30P140 U171 ( .A1(a[23]), .A2(n47), .A3(a[144]), .A4(n122), .Z(
        b[23]) );
  XOR4D1BWP30P140 U172 ( .A1(a[21]), .A2(n48), .A3(a[142]), .A4(n123), .Z(
        b[21]) );
  XOR4D1BWP30P140 U173 ( .A1(a[19]), .A2(n50), .A3(a[140]), .A4(n125), .Z(
        b[19]) );
  XOR4D1BWP30P140 U174 ( .A1(a[17]), .A2(n52), .A3(a[138]), .A4(n127), .Z(
        b[17]) );
  XOR4D1BWP30P140 U175 ( .A1(a[74]), .A2(a[200]), .A3(n29), .A4(n86), .Z(b[74]) );
  XOR4D1BWP30P140 U176 ( .A1(a[72]), .A2(a[198]), .A3(n30), .A4(n87), .Z(b[72]) );
  XOR4D1BWP30P140 U177 ( .A1(a[94]), .A2(a[220]), .A3(n18), .A4(n73), .Z(b[94]) );
  XOR4D1BWP30P140 U178 ( .A1(a[92]), .A2(a[218]), .A3(n19), .A4(n74), .Z(b[92]) );
  XOR4D1BWP30P140 U179 ( .A1(a[90]), .A2(a[216]), .A3(n20), .A4(n75), .Z(b[90]) );
  XOR4D1BWP30P140 U180 ( .A1(a[88]), .A2(a[214]), .A3(n21), .A4(n77), .Z(b[88]) );
  XOR4D1BWP30P140 U181 ( .A1(a[86]), .A2(a[212]), .A3(n22), .A4(n78), .Z(b[86]) );
  XOR4D1BWP30P140 U182 ( .A1(a[84]), .A2(a[210]), .A3(n23), .A4(n79), .Z(b[84]) );
  XOR4D1BWP30P140 U183 ( .A1(a[82]), .A2(a[208]), .A3(n24), .A4(n80), .Z(b[82]) );
  XOR4D1BWP30P140 U184 ( .A1(a[80]), .A2(a[206]), .A3(n25), .A4(n81), .Z(b[80]) );
  XOR4D1BWP30P140 U185 ( .A1(a[78]), .A2(a[204]), .A3(n26), .A4(n84), .Z(b[78]) );
  XOR4D1BWP30P140 U186 ( .A1(a[76]), .A2(a[202]), .A3(n27), .A4(n85), .Z(b[76]) );
  XOR4D1BWP30P140 U187 ( .A1(a[70]), .A2(a[196]), .A3(n31), .A4(n88), .Z(b[70]) );
  XOR4D1BWP30P140 U188 ( .A1(n67), .A2(n68), .A3(a[9]), .A4(a[137]), .Z(b[9])
         );
  XOR4D1BWP30P140 U189 ( .A1(n67), .A2(n76), .A3(a[8]), .A4(a[134]), .Z(b[8])
         );
  XOR4D1BWP30P140 U190 ( .A1(a[62]), .A2(n32), .A3(a[183]), .A4(n94), .Z(b[62]) );
  XOR4D1BWP30P140 U191 ( .A1(a[60]), .A2(n32), .A3(a[181]), .A4(n96), .Z(b[60]) );
  XOR4D1BWP30P140 U192 ( .A1(a[54]), .A2(n33), .A3(a[175]), .A4(n101), .Z(
        b[54]) );
  XOR4D1BWP30P140 U193 ( .A1(a[42]), .A2(n40), .A3(a[163]), .A4(n109), .Z(
        b[42]) );
  XOR4D1BWP30P140 U194 ( .A1(a[40]), .A2(n41), .A3(a[161]), .A4(n110), .Z(
        b[40]) );
  XOR4D1BWP30P140 U195 ( .A1(n82), .A2(n83), .A3(a[7]), .A4(a[135]), .Z(b[7])
         );
  XOR4D1BWP30P140 U196 ( .A1(a[36]), .A2(a[162]), .A3(n44), .A4(n113), .Z(
        b[36]) );
  XOR4D1BWP30P140 U197 ( .A1(a[34]), .A2(a[160]), .A3(n45), .A4(n114), .Z(
        b[34]) );
  XOR4D1BWP30P140 U198 ( .A1(a[52]), .A2(n34), .A3(a[173]), .A4(n102), .Z(
        b[52]) );
  XOR4D1BWP30P140 U199 ( .A1(a[50]), .A2(n35), .A3(a[171]), .A4(n103), .Z(
        b[50]) );
  XOR4D1BWP30P140 U200 ( .A1(a[48]), .A2(n36), .A3(a[169]), .A4(n105), .Z(
        b[48]) );
  XOR4D1BWP30P140 U201 ( .A1(a[46]), .A2(n37), .A3(a[167]), .A4(n106), .Z(
        b[46]) );
  XOR4D1BWP30P140 U202 ( .A1(a[15]), .A2(n53), .A3(a[136]), .A4(n128), .Z(
        b[15]) );
  XOR4D1BWP30P140 U203 ( .A1(a[44]), .A2(a[172]), .A3(n42), .A4(n108), .Z(
        b[44]) );
  XOR4D1BWP30P140 U204 ( .A1(n104), .A2(n135), .A3(a[139]), .A4(a[11]), .Z(
        b[11]) );
  XOR4D1BWP30P140 U205 ( .A1(a[32]), .A2(a[158]), .A3(n46), .A4(n115), .Z(
        b[32]) );
  XOR4D1BWP30P140 U206 ( .A1(a[30]), .A2(a[156]), .A3(n47), .A4(n116), .Z(
        b[30]) );
  XOR4D1BWP30P140 U207 ( .A1(a[28]), .A2(a[154]), .A3(n48), .A4(n119), .Z(
        b[28]) );
  XOR4D1BWP30P140 U208 ( .A1(a[26]), .A2(a[152]), .A3(n50), .A4(n120), .Z(
        b[26]) );
  XOR4D1BWP30P140 U209 ( .A1(a[24]), .A2(a[150]), .A3(n52), .A4(n121), .Z(
        b[24]) );
  XOR4D1BWP30P140 U210 ( .A1(a[22]), .A2(a[148]), .A3(n53), .A4(n122), .Z(
        b[22]) );
  XOR4D1BWP30P140 U211 ( .A1(n132), .A2(a[125]), .A3(a[251]), .A4(a[246]), .Z(
        b[125]) );
  XOR2UD1BWP30P140 U212 ( .A1(a[253]), .A2(a[252]), .Z(n132) );
  XOR4D1BWP30P140 U213 ( .A1(n97), .A2(n135), .A3(a[136]), .A4(a[10]), .Z(
        b[10]) );
  XOR4D1BWP30P140 U214 ( .A1(n97), .A2(n104), .A3(a[4]), .A4(n68), .Z(b[4]) );
  XOR4D1BWP30P140 U215 ( .A1(a[242]), .A2(a[116]), .A3(n7), .A4(n137), .Z(
        b[116]) );
  XOR4D1BWP30P140 U216 ( .A1(a[141]), .A2(a[13]), .A3(a[134]), .A4(n130), .Z(
        b[13]) );
  XOR4D1BWP30P140 U217 ( .A1(a[238]), .A2(a[112]), .A3(n9), .A4(n139), .Z(
        b[112]) );
  XOR4D1BWP30P140 U218 ( .A1(a[236]), .A2(a[110]), .A3(n10), .A4(n140), .Z(
        b[110]) );
  XOR4D1BWP30P140 U219 ( .A1(a[234]), .A2(a[108]), .A3(n11), .A4(n141), .Z(
        b[108]) );
  XOR4D1BWP30P140 U220 ( .A1(a[232]), .A2(a[106]), .A3(n12), .A4(n142), .Z(
        b[106]) );
  XOR4D1BWP30P140 U221 ( .A1(a[230]), .A2(a[104]), .A3(n14), .A4(n143), .Z(
        b[104]) );
  XOR4D1BWP30P140 U222 ( .A1(a[228]), .A2(a[102]), .A3(n16), .A4(n144), .Z(
        b[102]) );
  XOR4D1BWP30P140 U223 ( .A1(a[226]), .A2(a[100]), .A3(n17), .A4(n145), .Z(
        b[100]) );
  XOR4D1BWP30P140 U224 ( .A1(a[248]), .A2(a[120]), .A3(n5), .A4(n134), .Z(
        b[120]) );
  XOR4D1BWP30P140 U225 ( .A1(a[240]), .A2(a[114]), .A3(n8), .A4(n138), .Z(
        b[114]) );
  INVD1BWP30P140 U226 ( .I(a[172]), .ZN(n39) );
  INVD1BWP30P140 U227 ( .I(a[213]), .ZN(n19) );
  INVD1BWP30P140 U228 ( .I(a[207]), .ZN(n22) );
  INVD1BWP30P140 U229 ( .I(a[193]), .ZN(n30) );
  INVD1BWP30P140 U230 ( .I(a[205]), .ZN(n23) );
  INVD1BWP30P140 U231 ( .I(a[203]), .ZN(n24) );
  INVD1BWP30P140 U232 ( .I(a[201]), .ZN(n25) );
  INVD1BWP30P140 U233 ( .I(a[199]), .ZN(n26) );
  INVD1BWP30P140 U234 ( .I(a[197]), .ZN(n27) );
  INVD1BWP30P140 U235 ( .I(a[215]), .ZN(n18) );
  INVD1BWP30P140 U236 ( .I(a[211]), .ZN(n20) );
  INVD1BWP30P140 U237 ( .I(a[209]), .ZN(n21) );
  INVD1BWP30P140 U238 ( .I(a[221]), .ZN(n17) );
  INVD1BWP30P140 U239 ( .I(a[191]), .ZN(n31) );
  INVD1BWP30P140 U240 ( .I(a[188]), .ZN(n32) );
  INVD1BWP30P140 U241 ( .I(a[243]), .ZN(n4) );
  INVD1BWP30P140 U242 ( .I(a[241]), .ZN(n5) );
  INVD1BWP30P140 U243 ( .I(a[155]), .ZN(n45) );
  INVD1BWP30P140 U244 ( .I(a[153]), .ZN(n46) );
  INVD1BWP30P140 U245 ( .I(a[149]), .ZN(n48) );
  INVD1BWP30P140 U246 ( .I(a[143]), .ZN(n53) );
  INVD1BWP30P140 U247 ( .I(a[157]), .ZN(n44) );
  INVD1BWP30P140 U248 ( .I(a[151]), .ZN(n47) );
  INVD1BWP30P140 U249 ( .I(a[147]), .ZN(n50) );
  INVD1BWP30P140 U250 ( .I(a[145]), .ZN(n52) );
  INVD1BWP30P140 U251 ( .I(a[195]), .ZN(n29) );
  INVD1BWP30P140 U252 ( .I(a[165]), .ZN(n42) );
  XNR3UD1BWP30P140 U253 ( .A1(a[130]), .A2(a[129]), .A3(n118), .ZN(n111) );
  XOR3UD1BWP30P140 U254 ( .A1(a[248]), .A2(a[127]), .A3(n98), .Z(b[127]) );
  XNR3UD1BWP30P140 U255 ( .A1(a[2]), .A2(n111), .A3(n117), .ZN(b[2]) );
  XNR3UD1BWP30P140 U256 ( .A1(a[1]), .A2(n76), .A3(n117), .ZN(b[1]) );
  XNR3UD1BWP30P140 U257 ( .A1(a[6]), .A2(n82), .A3(n89), .ZN(b[6]) );
  XOR3UD1BWP30P140 U258 ( .A1(a[3]), .A2(n97), .A3(n111), .Z(b[3]) );
  XOR3UD1BWP30P140 U259 ( .A1(a[12]), .A2(n130), .A3(n131), .Z(b[12]) );
  XOR3UD1BWP30P140 U260 ( .A1(a[254]), .A2(a[138]), .A3(a[133]), .Z(n131) );
  INVD1BWP30P140 U261 ( .I(n129), .ZN(b_14_) );
  XOR4D1BWP30P140 U262 ( .A1(a[14]), .A2(a[140]), .A3(a[135]), .A4(n128), .Z(
        n129) );
  INVD1BWP30P140 U263 ( .I(n124), .ZN(b_20_) );
  XOR4D1BWP30P140 U264 ( .A1(a[20]), .A2(a[146]), .A3(a[141]), .A4(n123), .Z(
        n124) );
  INVD1BWP30P140 U265 ( .I(n126), .ZN(b_18_) );
  XOR4D1BWP30P140 U266 ( .A1(a[18]), .A2(a[144]), .A3(a[139]), .A4(n125), .Z(
        n126) );
endmodule
