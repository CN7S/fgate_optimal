module os_128bit_0 ( z0, z1, z2, y, C_g1, rst_n );
input [126:0] z0;
input [126:0] z1;
input [126:0] z2;
output [254:0] y;
input [21:0] C_g1;
input rst_n;
wire [126:0] _z0;
wire [126:0] _z1;
wire [126:0] _z2;
wire [254:0] _y;
wire [21:0] _C_g1;
wire _rst_n;
assign _y[0] = z0[0];
assign _z0[126:1] = z0[126:1];
assign _z1 = z1;
assign _z2[125:0] = z2[125:0];
assign _y[254] = z2[126];
assign y = _y;
assign _C_g1 = C_g1;
assign _rst_n = rst_n;
XOR3UD1BWP30P140 U0 ( .A1( _y[0] ), .A2( _z1[0] ), .A3( _z2[0] ), .Z( _y[1] ) );
XOR3UD1BWP30P140 U1 ( .A1( _z0[1] ), .A2( _z1[1] ), .A3( _z2[1] ), .Z( _y[3] ) );
XOR3UD1BWP30P140 U2 ( .A1( _z0[2] ), .A2( _z1[2] ), .A3( _z2[2] ), .Z( _y[5] ) );
XOR3UD1BWP30P140 U3 ( .A1( _z0[3] ), .A2( _z1[3] ), .A3( _z2[3] ), .Z( _y[7] ) );
XOR3UD1BWP30P140 U4 ( .A1( _z0[4] ), .A2( _z1[4] ), .A3( _z2[4] ), .Z( _y[9] ) );
XOR3UD1BWP30P140 U5 ( .A1( _z0[5] ), .A2( _z1[5] ), .A3( _z2[5] ), .Z( _y[11] ) );
XOR3UD1BWP30P140 U6 ( .A1( _z0[6] ), .A2( _z1[6] ), .A3( _z2[6] ), .Z( _y[13] ) );
XOR3UD1BWP30P140 U7 ( .A1( _z0[7] ), .A2( _z1[7] ), .A3( _z2[7] ), .Z( _y[15] ) );
XOR3UD1BWP30P140 U8 ( .A1( _z0[8] ), .A2( _z1[8] ), .A3( _z2[8] ), .Z( _y[17] ) );
XOR3UD1BWP30P140 U9 ( .A1( _z0[9] ), .A2( _z1[9] ), .A3( _z2[9] ), .Z( _y[19] ) );
XOR3UD1BWP30P140 U10 ( .A1( _z0[10] ), .A2( _z1[10] ), .A3( _z2[10] ), .Z( _y[21] ) );
XOR3UD1BWP30P140 U11 ( .A1( _z0[11] ), .A2( _z1[11] ), .A3( _z2[11] ), .Z( _y[23] ) );
XOR3UD1BWP30P140 U12 ( .A1( _z0[12] ), .A2( _z1[12] ), .A3( _z2[12] ), .Z( _y[25] ) );
XOR3UD1BWP30P140 U13 ( .A1( _z0[13] ), .A2( _z1[13] ), .A3( _z2[13] ), .Z( _y[27] ) );
XOR3UD1BWP30P140 U14 ( .A1( _z0[14] ), .A2( _z1[14] ), .A3( _z2[14] ), .Z( _y[29] ) );
XOR3UD1BWP30P140 U15 ( .A1( _z0[15] ), .A2( _z1[15] ), .A3( _z2[15] ), .Z( _y[31] ) );
XOR3UD1BWP30P140 U16 ( .A1( _z0[16] ), .A2( _z1[16] ), .A3( _z2[16] ), .Z( _y[33] ) );
XOR3UD1BWP30P140 U17 ( .A1( _z0[17] ), .A2( _z1[17] ), .A3( _z2[17] ), .Z( _y[35] ) );
XOR3UD1BWP30P140 U18 ( .A1( _z0[18] ), .A2( _z1[18] ), .A3( _z2[18] ), .Z( _y[37] ) );
XOR3UD1BWP30P140 U19 ( .A1( _z0[19] ), .A2( _z1[19] ), .A3( _z2[19] ), .Z( _y[39] ) );
XOR3UD1BWP30P140 U20 ( .A1( _z0[20] ), .A2( _z1[20] ), .A3( _z2[20] ), .Z( _y[41] ) );
XOR3UD1BWP30P140 U21 ( .A1( _z0[21] ), .A2( _z1[21] ), .A3( _z2[21] ), .Z( _y[43] ) );
XOR3UD1BWP30P140 U22 ( .A1( _z0[22] ), .A2( _z1[22] ), .A3( _z2[22] ), .Z( _y[45] ) );
XOR3UD1BWP30P140 U23 ( .A1( _z0[23] ), .A2( _z1[23] ), .A3( _z2[23] ), .Z( _y[47] ) );
XOR3UD1BWP30P140 U24 ( .A1( _z0[24] ), .A2( _z1[24] ), .A3( _z2[24] ), .Z( _y[49] ) );
XOR3UD1BWP30P140 U25 ( .A1( _z0[25] ), .A2( _z1[25] ), .A3( _z2[25] ), .Z( _y[51] ) );
XOR3UD1BWP30P140 U26 ( .A1( _z0[26] ), .A2( _z1[26] ), .A3( _z2[26] ), .Z( _y[53] ) );
XOR3UD1BWP30P140 U27 ( .A1( _z0[27] ), .A2( _z1[27] ), .A3( _z2[27] ), .Z( _y[55] ) );
XOR3UD1BWP30P140 U28 ( .A1( _z0[28] ), .A2( _z1[28] ), .A3( _z2[28] ), .Z( _y[57] ) );
XOR3UD1BWP30P140 U29 ( .A1( _z0[29] ), .A2( _z1[29] ), .A3( _z2[29] ), .Z( _y[59] ) );
XOR3UD1BWP30P140 U30 ( .A1( _z0[30] ), .A2( _z1[30] ), .A3( _z2[30] ), .Z( _y[61] ) );
XOR3UD1BWP30P140 U31 ( .A1( _z0[31] ), .A2( _z1[31] ), .A3( _z2[31] ), .Z( _y[63] ) );
XOR3UD1BWP30P140 U32 ( .A1( _z0[32] ), .A2( _z1[32] ), .A3( _z2[32] ), .Z( _y[65] ) );
XOR3UD1BWP30P140 U33 ( .A1( _z0[33] ), .A2( _z1[33] ), .A3( _z2[33] ), .Z( _y[67] ) );
XOR3UD1BWP30P140 U34 ( .A1( _z0[34] ), .A2( _z1[34] ), .A3( _z2[34] ), .Z( _y[69] ) );
XOR3UD1BWP30P140 U35 ( .A1( _z0[35] ), .A2( _z1[35] ), .A3( _z2[35] ), .Z( _y[71] ) );
XOR3UD1BWP30P140 U36 ( .A1( _z0[36] ), .A2( _z1[36] ), .A3( _z2[36] ), .Z( _y[73] ) );
XOR3UD1BWP30P140 U37 ( .A1( _z0[37] ), .A2( _z1[37] ), .A3( _z2[37] ), .Z( _y[75] ) );
XOR3UD1BWP30P140 U38 ( .A1( _z0[38] ), .A2( _z1[38] ), .A3( _z2[38] ), .Z( _y[77] ) );
XOR3UD1BWP30P140 U39 ( .A1( _z0[39] ), .A2( _z1[39] ), .A3( _z2[39] ), .Z( _y[79] ) );
XOR3UD1BWP30P140 U40 ( .A1( _z0[40] ), .A2( _z1[40] ), .A3( _z2[40] ), .Z( _y[81] ) );
XOR3UD1BWP30P140 U41 ( .A1( _z0[41] ), .A2( _z1[41] ), .A3( _z2[41] ), .Z( _y[83] ) );
XOR3UD1BWP30P140 U42 ( .A1( _z0[42] ), .A2( _z1[42] ), .A3( _z2[42] ), .Z( _y[85] ) );
XOR3UD1BWP30P140 U43 ( .A1( _z0[43] ), .A2( _z1[43] ), .A3( _z2[43] ), .Z( _y[87] ) );
XOR3UD1BWP30P140 U44 ( .A1( _z0[44] ), .A2( _z1[44] ), .A3( _z2[44] ), .Z( _y[89] ) );
XOR3UD1BWP30P140 U45 ( .A1( _z0[45] ), .A2( _z1[45] ), .A3( _z2[45] ), .Z( _y[91] ) );
XOR3UD1BWP30P140 U46 ( .A1( _z0[46] ), .A2( _z1[46] ), .A3( _z2[46] ), .Z( _y[93] ) );
XOR3UD1BWP30P140 U47 ( .A1( _z0[47] ), .A2( _z1[47] ), .A3( _z2[47] ), .Z( _y[95] ) );
XOR3UD1BWP30P140 U48 ( .A1( _z0[48] ), .A2( _z1[48] ), .A3( _z2[48] ), .Z( _y[97] ) );
XOR3UD1BWP30P140 U49 ( .A1( _z0[49] ), .A2( _z1[49] ), .A3( _z2[49] ), .Z( _y[99] ) );
XOR3UD1BWP30P140 U50 ( .A1( _z0[50] ), .A2( _z1[50] ), .A3( _z2[50] ), .Z( _y[101] ) );
XOR3UD1BWP30P140 U51 ( .A1( _z0[51] ), .A2( _z1[51] ), .A3( _z2[51] ), .Z( _y[103] ) );
XOR3UD1BWP30P140 U52 ( .A1( _z0[52] ), .A2( _z1[52] ), .A3( _z2[52] ), .Z( _y[105] ) );
XOR3UD1BWP30P140 U53 ( .A1( _z0[53] ), .A2( _z1[53] ), .A3( _z2[53] ), .Z( _y[107] ) );
XOR3UD1BWP30P140 U54 ( .A1( _z0[54] ), .A2( _z1[54] ), .A3( _z2[54] ), .Z( _y[109] ) );
XOR3UD1BWP30P140 U55 ( .A1( _z0[55] ), .A2( _z1[55] ), .A3( _z2[55] ), .Z( _y[111] ) );
XOR3UD1BWP30P140 U56 ( .A1( _z0[56] ), .A2( _z1[56] ), .A3( _z2[56] ), .Z( _y[113] ) );
XOR3UD1BWP30P140 U57 ( .A1( _z0[57] ), .A2( _z1[57] ), .A3( _z2[57] ), .Z( _y[115] ) );
XOR3UD1BWP30P140 U58 ( .A1( _z0[58] ), .A2( _z1[58] ), .A3( _z2[58] ), .Z( _y[117] ) );
XOR3UD1BWP30P140 U59 ( .A1( _z0[59] ), .A2( _z1[59] ), .A3( _z2[59] ), .Z( _y[119] ) );
XOR3UD1BWP30P140 U60 ( .A1( _z0[60] ), .A2( _z1[60] ), .A3( _z2[60] ), .Z( _y[121] ) );
XOR3UD1BWP30P140 U61 ( .A1( _z0[61] ), .A2( _z1[61] ), .A3( _z2[61] ), .Z( _y[123] ) );
XOR3UD1BWP30P140 U62 ( .A1( _z0[62] ), .A2( _z1[62] ), .A3( _z2[62] ), .Z( _y[125] ) );
XOR3UD1BWP30P140 U63 ( .A1( _z0[63] ), .A2( _z1[63] ), .A3( _z2[63] ), .Z( _y[127] ) );
XOR3UD1BWP30P140 U64 ( .A1( _z0[64] ), .A2( _z1[64] ), .A3( _z2[64] ), .Z( _y[129] ) );
XOR3UD1BWP30P140 U65 ( .A1( _z0[65] ), .A2( _z1[65] ), .A3( _z2[65] ), .Z( _y[131] ) );
XOR3UD1BWP30P140 U66 ( .A1( _z0[66] ), .A2( _z1[66] ), .A3( _z2[66] ), .Z( _y[133] ) );
XOR3UD1BWP30P140 U67 ( .A1( _z0[67] ), .A2( _z1[67] ), .A3( _z2[67] ), .Z( _y[135] ) );
XOR3UD1BWP30P140 U68 ( .A1( _z0[68] ), .A2( _z1[68] ), .A3( _z2[68] ), .Z( _y[137] ) );
XOR3UD1BWP30P140 U69 ( .A1( _z0[69] ), .A2( _z1[69] ), .A3( _z2[69] ), .Z( _y[139] ) );
XOR3UD1BWP30P140 U70 ( .A1( _z0[70] ), .A2( _z1[70] ), .A3( _z2[70] ), .Z( _y[141] ) );
XOR3UD1BWP30P140 U71 ( .A1( _z0[71] ), .A2( _z1[71] ), .A3( _z2[71] ), .Z( _y[143] ) );
XOR3UD1BWP30P140 U72 ( .A1( _z0[72] ), .A2( _z1[72] ), .A3( _z2[72] ), .Z( _y[145] ) );
XOR3UD1BWP30P140 U73 ( .A1( _z0[73] ), .A2( _z1[73] ), .A3( _z2[73] ), .Z( _y[147] ) );
XOR3UD1BWP30P140 U74 ( .A1( _z0[74] ), .A2( _z1[74] ), .A3( _z2[74] ), .Z( _y[149] ) );
XOR3UD1BWP30P140 U75 ( .A1( _z0[75] ), .A2( _z1[75] ), .A3( _z2[75] ), .Z( _y[151] ) );
XOR3UD1BWP30P140 U76 ( .A1( _z0[76] ), .A2( _z1[76] ), .A3( _z2[76] ), .Z( _y[153] ) );
XOR3UD1BWP30P140 U77 ( .A1( _z0[77] ), .A2( _z1[77] ), .A3( _z2[77] ), .Z( _y[155] ) );
XOR3UD1BWP30P140 U78 ( .A1( _z0[78] ), .A2( _z1[78] ), .A3( _z2[78] ), .Z( _y[157] ) );
XOR3UD1BWP30P140 U79 ( .A1( _z0[79] ), .A2( _z1[79] ), .A3( _z2[79] ), .Z( _y[159] ) );
XOR3UD1BWP30P140 U80 ( .A1( _z0[80] ), .A2( _z1[80] ), .A3( _z2[80] ), .Z( _y[161] ) );
XOR3UD1BWP30P140 U81 ( .A1( _z0[81] ), .A2( _z1[81] ), .A3( _z2[81] ), .Z( _y[163] ) );
XOR3UD1BWP30P140 U82 ( .A1( _z0[82] ), .A2( _z1[82] ), .A3( _z2[82] ), .Z( _y[165] ) );
XOR3UD1BWP30P140 U83 ( .A1( _z0[83] ), .A2( _z1[83] ), .A3( _z2[83] ), .Z( _y[167] ) );
XOR3UD1BWP30P140 U84 ( .A1( _z0[84] ), .A2( _z1[84] ), .A3( _z2[84] ), .Z( _y[169] ) );
XOR3UD1BWP30P140 U85 ( .A1( _z0[85] ), .A2( _z1[85] ), .A3( _z2[85] ), .Z( _y[171] ) );
XOR3UD1BWP30P140 U86 ( .A1( _z0[86] ), .A2( _z1[86] ), .A3( _z2[86] ), .Z( _y[173] ) );
XOR3UD1BWP30P140 U87 ( .A1( _z0[87] ), .A2( _z1[87] ), .A3( _z2[87] ), .Z( _y[175] ) );
XOR3UD1BWP30P140 U88 ( .A1( _z0[88] ), .A2( _z1[88] ), .A3( _z2[88] ), .Z( _y[177] ) );
XOR3UD1BWP30P140 U89 ( .A1( _z0[89] ), .A2( _z1[89] ), .A3( _z2[89] ), .Z( _y[179] ) );
XOR3UD1BWP30P140 U90 ( .A1( _z0[90] ), .A2( _z1[90] ), .A3( _z2[90] ), .Z( _y[181] ) );
XOR3UD1BWP30P140 U91 ( .A1( _z0[91] ), .A2( _z1[91] ), .A3( _z2[91] ), .Z( _y[183] ) );
XOR3UD1BWP30P140 U92 ( .A1( _z0[92] ), .A2( _z1[92] ), .A3( _z2[92] ), .Z( _y[185] ) );
XOR3UD1BWP30P140 U93 ( .A1( _z0[93] ), .A2( _z1[93] ), .A3( _z2[93] ), .Z( _y[187] ) );
XOR3UD1BWP30P140 U94 ( .A1( _z0[94] ), .A2( _z1[94] ), .A3( _z2[94] ), .Z( _y[189] ) );
XOR3UD1BWP30P140 U95 ( .A1( _z0[95] ), .A2( _z1[95] ), .A3( _z2[95] ), .Z( _y[191] ) );
XOR3UD1BWP30P140 U96 ( .A1( _z0[96] ), .A2( _z1[96] ), .A3( _z2[96] ), .Z( _y[193] ) );
XOR3UD1BWP30P140 U97 ( .A1( _z0[97] ), .A2( _z1[97] ), .A3( _z2[97] ), .Z( _y[195] ) );
XOR3UD1BWP30P140 U98 ( .A1( _z0[98] ), .A2( _z1[98] ), .A3( _z2[98] ), .Z( _y[197] ) );
XOR3UD1BWP30P140 U99 ( .A1( _z0[99] ), .A2( _z1[99] ), .A3( _z2[99] ), .Z( _y[199] ) );
XOR3UD1BWP30P140 U100 ( .A1( _z0[100] ), .A2( _z1[100] ), .A3( _z2[100] ), .Z( _y[201] ) );
XOR3UD1BWP30P140 U101 ( .A1( _z0[101] ), .A2( _z1[101] ), .A3( _z2[101] ), .Z( _y[203] ) );
XOR3UD1BWP30P140 U102 ( .A1( _z0[102] ), .A2( _z1[102] ), .A3( _z2[102] ), .Z( _y[205] ) );
XOR3UD1BWP30P140 U103 ( .A1( _z0[103] ), .A2( _z1[103] ), .A3( _z2[103] ), .Z( _y[207] ) );
XOR3UD1BWP30P140 U104 ( .A1( _z0[104] ), .A2( _z1[104] ), .A3( _z2[104] ), .Z( _y[209] ) );
XOR3UD1BWP30P140 U105 ( .A1( _z0[105] ), .A2( _z1[105] ), .A3( _z2[105] ), .Z( _y[211] ) );
XOR3UD1BWP30P140 U106 ( .A1( _z0[106] ), .A2( _z1[106] ), .A3( _z2[106] ), .Z( _y[213] ) );
XOR3UD1BWP30P140 U107 ( .A1( _z0[107] ), .A2( _z1[107] ), .A3( _z2[107] ), .Z( _y[215] ) );
XOR3UD1BWP30P140 U108 ( .A1( _z0[108] ), .A2( _z1[108] ), .A3( _z2[108] ), .Z( _y[217] ) );
XOR3UD1BWP30P140 U109 ( .A1( _z0[109] ), .A2( _z1[109] ), .A3( _z2[109] ), .Z( _y[219] ) );
XOR3UD1BWP30P140 U110 ( .A1( _z0[110] ), .A2( _z1[110] ), .A3( _z2[110] ), .Z( _y[221] ) );
XOR3UD1BWP30P140 U111 ( .A1( _z0[111] ), .A2( _z1[111] ), .A3( _z2[111] ), .Z( _y[223] ) );
XOR3UD1BWP30P140 U112 ( .A1( _z0[112] ), .A2( _z1[112] ), .A3( _z2[112] ), .Z( _y[225] ) );
XOR3UD1BWP30P140 U113 ( .A1( _z0[113] ), .A2( _z1[113] ), .A3( _z2[113] ), .Z( _y[227] ) );
XOR3UD1BWP30P140 U114 ( .A1( _z0[114] ), .A2( _z1[114] ), .A3( _z2[114] ), .Z( _y[229] ) );
XOR3UD1BWP30P140 U115 ( .A1( _z0[115] ), .A2( _z1[115] ), .A3( _z2[115] ), .Z( _y[231] ) );
XOR3UD1BWP30P140 U116 ( .A1( _z0[116] ), .A2( _z1[116] ), .A3( _z2[116] ), .Z( _y[233] ) );
XOR3UD1BWP30P140 U117 ( .A1( _z0[117] ), .A2( _z1[117] ), .A3( _z2[117] ), .Z( _y[235] ) );
XOR3UD1BWP30P140 U118 ( .A1( _z0[118] ), .A2( _z1[118] ), .A3( _z2[118] ), .Z( _y[237] ) );
XOR3UD1BWP30P140 U119 ( .A1( _z0[119] ), .A2( _z1[119] ), .A3( _z2[119] ), .Z( _y[239] ) );
XOR3UD1BWP30P140 U120 ( .A1( _z0[120] ), .A2( _z1[120] ), .A3( _z2[120] ), .Z( _y[241] ) );
XOR3UD1BWP30P140 U121 ( .A1( _z0[121] ), .A2( _z1[121] ), .A3( _z2[121] ), .Z( _y[243] ) );
XOR3UD1BWP30P140 U122 ( .A1( _z0[122] ), .A2( _z1[122] ), .A3( _z2[122] ), .Z( _y[245] ) );
XOR3UD1BWP30P140 U123 ( .A1( _z0[123] ), .A2( _z1[123] ), .A3( _z2[123] ), .Z( _y[247] ) );
XOR3UD1BWP30P140 U124 ( .A1( _z0[124] ), .A2( _z1[124] ), .A3( _z2[124] ), .Z( _y[249] ) );
XOR3UD1BWP30P140 U125 ( .A1( _z0[125] ), .A2( _z1[125] ), .A3( _z2[125] ), .Z( _y[251] ) );
XOR3UD1BWP30P140 U126 ( .A1( _z0[126] ), .A2( _z1[126] ), .A3( _y[254] ), .Z( _y[253] ) );
XOR2UD1BWP30P140 U127 ( .A1( _z0[1] ), .A2( _z2[0] ), .Z( _y[2] ) );
XOR2UD1BWP30P140 U128 ( .A1( _z0[2] ), .A2( _z2[1] ), .Z( _y[4] ) );
XOR2UD1BWP30P140 U129 ( .A1( _z0[3] ), .A2( _z2[2] ), .Z( _y[6] ) );
XOR2UD1BWP30P140 U130 ( .A1( _z0[4] ), .A2( _z2[3] ), .Z( _y[8] ) );
XOR2UD1BWP30P140 U131 ( .A1( _z0[5] ), .A2( _z2[4] ), .Z( _y[10] ) );
XOR2UD1BWP30P140 U132 ( .A1( _z0[6] ), .A2( _z2[5] ), .Z( _y[12] ) );
XOR2UD1BWP30P140 U133 ( .A1( _z0[7] ), .A2( _z2[6] ), .Z( _y[14] ) );
XOR2UD1BWP30P140 U134 ( .A1( _z0[8] ), .A2( _z2[7] ), .Z( _y[16] ) );
XOR2UD1BWP30P140 U135 ( .A1( _z0[9] ), .A2( _z2[8] ), .Z( _y[18] ) );
XOR2UD1BWP30P140 U136 ( .A1( _z0[10] ), .A2( _z2[9] ), .Z( _y[20] ) );
XOR2UD1BWP30P140 U137 ( .A1( _z0[11] ), .A2( _z2[10] ), .Z( _y[22] ) );
XOR2UD1BWP30P140 U138 ( .A1( _z0[12] ), .A2( _z2[11] ), .Z( _y[24] ) );
XOR2UD1BWP30P140 U139 ( .A1( _z0[13] ), .A2( _z2[12] ), .Z( _y[26] ) );
XOR2UD1BWP30P140 U140 ( .A1( _z0[14] ), .A2( _z2[13] ), .Z( _y[28] ) );
XOR2UD1BWP30P140 U141 ( .A1( _z0[15] ), .A2( _z2[14] ), .Z( _y[30] ) );
XOR2UD1BWP30P140 U142 ( .A1( _z0[16] ), .A2( _z2[15] ), .Z( _y[32] ) );
XOR2UD1BWP30P140 U143 ( .A1( _z0[17] ), .A2( _z2[16] ), .Z( _y[34] ) );
XOR2UD1BWP30P140 U144 ( .A1( _z0[18] ), .A2( _z2[17] ), .Z( _y[36] ) );
XOR2UD1BWP30P140 U145 ( .A1( _z0[19] ), .A2( _z2[18] ), .Z( _y[38] ) );
XOR2UD1BWP30P140 U146 ( .A1( _z0[20] ), .A2( _z2[19] ), .Z( _y[40] ) );
XOR2UD1BWP30P140 U147 ( .A1( _z0[21] ), .A2( _z2[20] ), .Z( _y[42] ) );
XOR2UD1BWP30P140 U148 ( .A1( _z0[22] ), .A2( _z2[21] ), .Z( _y[44] ) );
XOR2UD1BWP30P140 U149 ( .A1( _z0[23] ), .A2( _z2[22] ), .Z( _y[46] ) );
XOR2UD1BWP30P140 U150 ( .A1( _z0[24] ), .A2( _z2[23] ), .Z( _y[48] ) );
XOR2UD1BWP30P140 U151 ( .A1( _z0[25] ), .A2( _z2[24] ), .Z( _y[50] ) );
XOR2UD1BWP30P140 U152 ( .A1( _z0[26] ), .A2( _z2[25] ), .Z( _y[52] ) );
XOR2UD1BWP30P140 U153 ( .A1( _z0[27] ), .A2( _z2[26] ), .Z( _y[54] ) );
XOR2UD1BWP30P140 U154 ( .A1( _z0[28] ), .A2( _z2[27] ), .Z( _y[56] ) );
XOR2UD1BWP30P140 U155 ( .A1( _z0[29] ), .A2( _z2[28] ), .Z( _y[58] ) );
XOR2UD1BWP30P140 U156 ( .A1( _z0[30] ), .A2( _z2[29] ), .Z( _y[60] ) );
XOR2UD1BWP30P140 U157 ( .A1( _z0[31] ), .A2( _z2[30] ), .Z( _y[62] ) );
XOR2UD1BWP30P140 U158 ( .A1( _z0[32] ), .A2( _z2[31] ), .Z( _y[64] ) );
XOR2UD1BWP30P140 U159 ( .A1( _z0[33] ), .A2( _z2[32] ), .Z( _y[66] ) );
XOR2UD1BWP30P140 U160 ( .A1( _z0[34] ), .A2( _z2[33] ), .Z( _y[68] ) );
XOR2UD1BWP30P140 U161 ( .A1( _z0[35] ), .A2( _z2[34] ), .Z( _y[70] ) );
XOR2UD1BWP30P140 U162 ( .A1( _z0[36] ), .A2( _z2[35] ), .Z( _y[72] ) );
XOR2UD1BWP30P140 U163 ( .A1( _z0[37] ), .A2( _z2[36] ), .Z( _y[74] ) );
XOR2UD1BWP30P140 U164 ( .A1( _z0[38] ), .A2( _z2[37] ), .Z( _y[76] ) );
XOR2UD1BWP30P140 U165 ( .A1( _z0[39] ), .A2( _z2[38] ), .Z( _y[78] ) );
XOR2UD1BWP30P140 U166 ( .A1( _z0[40] ), .A2( _z2[39] ), .Z( _y[80] ) );
XOR2UD1BWP30P140 U167 ( .A1( _z0[41] ), .A2( _z2[40] ), .Z( _y[82] ) );
XOR2UD1BWP30P140 U168 ( .A1( _z0[42] ), .A2( _z2[41] ), .Z( _y[84] ) );
XOR2UD1BWP30P140 U169 ( .A1( _z0[43] ), .A2( _z2[42] ), .Z( _y[86] ) );
XOR2UD1BWP30P140 U170 ( .A1( _z0[44] ), .A2( _z2[43] ), .Z( _y[88] ) );
XOR2UD1BWP30P140 U171 ( .A1( _z0[45] ), .A2( _z2[44] ), .Z( _y[90] ) );
XOR2UD1BWP30P140 U172 ( .A1( _z0[46] ), .A2( _z2[45] ), .Z( _y[92] ) );
XOR2UD1BWP30P140 U173 ( .A1( _z0[47] ), .A2( _z2[46] ), .Z( _y[94] ) );
XOR2UD1BWP30P140 U174 ( .A1( _z0[48] ), .A2( _z2[47] ), .Z( _y[96] ) );
XOR2UD1BWP30P140 U175 ( .A1( _z0[49] ), .A2( _z2[48] ), .Z( _y[98] ) );
XOR2UD1BWP30P140 U176 ( .A1( _z0[50] ), .A2( _z2[49] ), .Z( _y[100] ) );
XOR2UD1BWP30P140 U177 ( .A1( _z0[51] ), .A2( _z2[50] ), .Z( _y[102] ) );
XOR2UD1BWP30P140 U178 ( .A1( _z0[52] ), .A2( _z2[51] ), .Z( _y[104] ) );
XOR2UD1BWP30P140 U179 ( .A1( _z0[53] ), .A2( _z2[52] ), .Z( _y[106] ) );
XOR2UD1BWP30P140 U180 ( .A1( _z0[54] ), .A2( _z2[53] ), .Z( _y[108] ) );
XOR2UD1BWP30P140 U181 ( .A1( _z0[55] ), .A2( _z2[54] ), .Z( _y[110] ) );
XOR2UD1BWP30P140 U182 ( .A1( _z0[56] ), .A2( _z2[55] ), .Z( _y[112] ) );
XOR2UD1BWP30P140 U183 ( .A1( _z0[57] ), .A2( _z2[56] ), .Z( _y[114] ) );
XOR2UD1BWP30P140 U184 ( .A1( _z0[58] ), .A2( _z2[57] ), .Z( _y[116] ) );
XOR2UD1BWP30P140 U185 ( .A1( _z0[59] ), .A2( _z2[58] ), .Z( _y[118] ) );
XOR2UD1BWP30P140 U186 ( .A1( _z0[60] ), .A2( _z2[59] ), .Z( _y[120] ) );
XOR2UD1BWP30P140 U187 ( .A1( _z0[61] ), .A2( _z2[60] ), .Z( _y[122] ) );
XOR2UD1BWP30P140 U188 ( .A1( _z0[62] ), .A2( _z2[61] ), .Z( _y[124] ) );
XOR2UD1BWP30P140 U189 ( .A1( _z0[63] ), .A2( _z2[62] ), .Z( _y[126] ) );
XOR2UD1BWP30P140 U190 ( .A1( _z0[64] ), .A2( _z2[63] ), .Z( _y[128] ) );
XOR2UD1BWP30P140 U191 ( .A1( _z0[65] ), .A2( _z2[64] ), .Z( _y[130] ) );
XOR2UD1BWP30P140 U192 ( .A1( _z0[66] ), .A2( _z2[65] ), .Z( _y[132] ) );
XOR2UD1BWP30P140 U193 ( .A1( _z0[67] ), .A2( _z2[66] ), .Z( _y[134] ) );
XOR2UD1BWP30P140 U194 ( .A1( _z0[68] ), .A2( _z2[67] ), .Z( _y[136] ) );
XOR2UD1BWP30P140 U195 ( .A1( _z0[69] ), .A2( _z2[68] ), .Z( _y[138] ) );
XOR2UD1BWP30P140 U196 ( .A1( _z0[70] ), .A2( _z2[69] ), .Z( _y[140] ) );
XOR2UD1BWP30P140 U197 ( .A1( _z0[71] ), .A2( _z2[70] ), .Z( _y[142] ) );
XOR2UD1BWP30P140 U198 ( .A1( _z0[72] ), .A2( _z2[71] ), .Z( _y[144] ) );
XOR2UD1BWP30P140 U199 ( .A1( _z0[73] ), .A2( _z2[72] ), .Z( _y[146] ) );
XOR2UD1BWP30P140 U200 ( .A1( _z0[74] ), .A2( _z2[73] ), .Z( _y[148] ) );
XOR2UD1BWP30P140 U201 ( .A1( _z0[75] ), .A2( _z2[74] ), .Z( _y[150] ) );
XOR2UD1BWP30P140 U202 ( .A1( _z0[76] ), .A2( _z2[75] ), .Z( _y[152] ) );
XOR2UD1BWP30P140 U203 ( .A1( _z0[77] ), .A2( _z2[76] ), .Z( _y[154] ) );
XOR2UD1BWP30P140 U204 ( .A1( _z0[78] ), .A2( _z2[77] ), .Z( _y[156] ) );
XOR2UD1BWP30P140 U205 ( .A1( _z0[79] ), .A2( _z2[78] ), .Z( _y[158] ) );
XOR2UD1BWP30P140 U206 ( .A1( _z0[80] ), .A2( _z2[79] ), .Z( _y[160] ) );
XOR2UD1BWP30P140 U207 ( .A1( _z0[81] ), .A2( _z2[80] ), .Z( _y[162] ) );
XOR2UD1BWP30P140 U208 ( .A1( _z0[82] ), .A2( _z2[81] ), .Z( _y[164] ) );
XOR2UD1BWP30P140 U209 ( .A1( _z0[83] ), .A2( _z2[82] ), .Z( _y[166] ) );
XOR2UD1BWP30P140 U210 ( .A1( _z0[84] ), .A2( _z2[83] ), .Z( _y[168] ) );
XOR2UD1BWP30P140 U211 ( .A1( _z0[85] ), .A2( _z2[84] ), .Z( _y[170] ) );
XOR2UD1BWP30P140 U212 ( .A1( _z0[86] ), .A2( _z2[85] ), .Z( _y[172] ) );
XOR2UD1BWP30P140 U213 ( .A1( _z0[87] ), .A2( _z2[86] ), .Z( _y[174] ) );
XOR2UD1BWP30P140 U214 ( .A1( _z0[88] ), .A2( _z2[87] ), .Z( _y[176] ) );
XOR2UD1BWP30P140 U215 ( .A1( _z0[89] ), .A2( _z2[88] ), .Z( _y[178] ) );
XOR2UD1BWP30P140 U216 ( .A1( _z0[90] ), .A2( _z2[89] ), .Z( _y[180] ) );
XOR2UD1BWP30P140 U217 ( .A1( _z0[91] ), .A2( _z2[90] ), .Z( _y[182] ) );
XOR2UD1BWP30P140 U218 ( .A1( _z0[92] ), .A2( _z2[91] ), .Z( _y[184] ) );
XOR2UD1BWP30P140 U219 ( .A1( _z0[93] ), .A2( _z2[92] ), .Z( _y[186] ) );
XOR2UD1BWP30P140 U220 ( .A1( _z0[94] ), .A2( _z2[93] ), .Z( _y[188] ) );
XOR2UD1BWP30P140 U221 ( .A1( _z0[95] ), .A2( _z2[94] ), .Z( _y[190] ) );
XOR2UD1BWP30P140 U222 ( .A1( _z0[96] ), .A2( _z2[95] ), .Z( _y[192] ) );
XOR2UD1BWP30P140 U223 ( .A1( _z0[97] ), .A2( _z2[96] ), .Z( _y[194] ) );
XOR2UD1BWP30P140 U224 ( .A1( _z0[98] ), .A2( _z2[97] ), .Z( _y[196] ) );
XOR2UD1BWP30P140 U225 ( .A1( _z0[99] ), .A2( _z2[98] ), .Z( _y[198] ) );
XOR2UD1BWP30P140 U226 ( .A1( _z0[100] ), .A2( _z2[99] ), .Z( _y[200] ) );
XOR2UD1BWP30P140 U227 ( .A1( _z0[101] ), .A2( _z2[100] ), .Z( _y[202] ) );
XOR2UD1BWP30P140 U228 ( .A1( _z0[102] ), .A2( _z2[101] ), .Z( _y[204] ) );
XOR2UD1BWP30P140 U229 ( .A1( _z0[103] ), .A2( _z2[102] ), .Z( _y[206] ) );
XOR2UD1BWP30P140 U230 ( .A1( _z0[104] ), .A2( _z2[103] ), .Z( _y[208] ) );
XOR2UD1BWP30P140 U231 ( .A1( _z0[105] ), .A2( _z2[104] ), .Z( _y[210] ) );
XOR2UD1BWP30P140 U232 ( .A1( _z0[106] ), .A2( _z2[105] ), .Z( _y[212] ) );
XOR2UD1BWP30P140 U233 ( .A1( _z0[107] ), .A2( _z2[106] ), .Z( _y[214] ) );
XOR2UD1BWP30P140 U234 ( .A1( _z0[108] ), .A2( _z2[107] ), .Z( _y[216] ) );
XOR2UD1BWP30P140 U235 ( .A1( _z0[109] ), .A2( _z2[108] ), .Z( _y[218] ) );
XOR2UD1BWP30P140 U236 ( .A1( _z0[110] ), .A2( _z2[109] ), .Z( _y[220] ) );
XOR2UD1BWP30P140 U237 ( .A1( _z0[111] ), .A2( _z2[110] ), .Z( _y[222] ) );
XOR2UD1BWP30P140 U238 ( .A1( _z0[112] ), .A2( _z2[111] ), .Z( _y[224] ) );
XOR2UD1BWP30P140 U239 ( .A1( _z0[113] ), .A2( _z2[112] ), .Z( _y[226] ) );
XOR2UD1BWP30P140 U240 ( .A1( _z0[114] ), .A2( _z2[113] ), .Z( _y[228] ) );
XOR2UD1BWP30P140 U241 ( .A1( _z0[115] ), .A2( _z2[114] ), .Z( _y[230] ) );
XOR2UD1BWP30P140 U242 ( .A1( _z0[116] ), .A2( _z2[115] ), .Z( _y[232] ) );
XOR2UD1BWP30P140 U243 ( .A1( _z0[117] ), .A2( _z2[116] ), .Z( _y[234] ) );
XOR2UD1BWP30P140 U244 ( .A1( _z0[118] ), .A2( _z2[117] ), .Z( _y[236] ) );
XOR2UD1BWP30P140 U245 ( .A1( _z0[119] ), .A2( _z2[118] ), .Z( _y[238] ) );
XOR2UD1BWP30P140 U246 ( .A1( _z0[120] ), .A2( _z2[119] ), .Z( _y[240] ) );
XOR2UD1BWP30P140 U247 ( .A1( _z0[121] ), .A2( _z2[120] ), .Z( _y[242] ) );
XOR2UD1BWP30P140 U248 ( .A1( _z0[122] ), .A2( _z2[121] ), .Z( _y[244] ) );
XOR2UD1BWP30P140 U249 ( .A1( _z0[123] ), .A2( _z2[122] ), .Z( _y[246] ) );
XOR2UD1BWP30P140 U250 ( .A1( _z0[124] ), .A2( _z2[123] ), .Z( _y[248] ) );
XOR2UD1BWP30P140 U251 ( .A1( _z0[125] ), .A2( _z2[124] ), .Z( _y[250] ) );
XOR2UD1BWP30P140 U252 ( .A1( _z0[126] ), .A2( _z2[125] ), .Z( _y[252] ) );
endmodule
